
module openMSP430(aclk, aclk_en, dbg_freeze, dbg_i2c_sda_out, dbg_uart_txd, dco_enable, dco_wkup, dmem_addr_0_, dmem_addr_1_, dmem_addr_2_, dmem_addr_3_, dmem_addr_4_, dmem_addr_5_, dmem_addr_6_, dmem_addr_7_, dmem_addr_8_, dmem_addr_9_, dmem_addr_10_, dmem_addr_11_, dmem_addr_12_, dmem_cen, dmem_din_0_, dmem_din_1_, dmem_din_2_, dmem_din_3_, dmem_din_4_, dmem_din_5_, dmem_din_6_, dmem_din_7_, dmem_din_8_, dmem_din_9_, dmem_din_10_, dmem_din_11_, dmem_din_12_, dmem_din_13_, dmem_din_14_, dmem_din_15_, dmem_wen_0_, dmem_wen_1_, irq_acc_0_, irq_acc_1_, irq_acc_2_, irq_acc_3_, irq_acc_4_, irq_acc_5_, irq_acc_6_, irq_acc_7_, irq_acc_8_, irq_acc_9_, irq_acc_10_, irq_acc_11_, irq_acc_12_, irq_acc_13_, lfxt_enable, lfxt_wkup, mclk, dma_dout_0_, dma_dout_1_, dma_dout_2_, dma_dout_3_, dma_dout_4_, dma_dout_5_, dma_dout_6_, dma_dout_7_, dma_dout_8_, dma_dout_9_, dma_dout_10_, dma_dout_11_, dma_dout_12_, dma_dout_13_, dma_dout_14_, dma_dout_15_, dma_ready, dma_resp, per_addr_0_, per_addr_1_, per_addr_2_, per_addr_3_, per_addr_4_, per_addr_5_, per_addr_6_, per_addr_7_, per_addr_8_, per_addr_9_, per_addr_10_, per_addr_11_, per_addr_12_, per_addr_13_, per_din_0_, per_din_1_, per_din_2_, per_din_3_, per_din_4_, per_din_5_, per_din_6_, per_din_7_, per_din_8_, per_din_9_, per_din_10_, per_din_11_, per_din_12_, per_din_13_, per_din_14_, per_din_15_, per_en, per_we_0_, per_we_1_, pmem_addr_0_, pmem_addr_1_, pmem_addr_2_, pmem_addr_3_, pmem_addr_4_, pmem_addr_5_, pmem_addr_6_, pmem_addr_7_, pmem_addr_8_, pmem_addr_9_, pmem_addr_10_, pmem_addr_11_, pmem_addr_12_, pmem_addr_13_, pmem_cen, pmem_din_0_, pmem_din_1_, pmem_din_2_, pmem_din_3_, pmem_din_4_, pmem_din_5_, pmem_din_6_, pmem_din_7_, pmem_din_8_, pmem_din_9_, pmem_din_10_, pmem_din_11_, pmem_din_12_, pmem_din_13_, pmem_din_14_, pmem_din_15_, pmem_wen_0_, pmem_wen_1_, puc_rst, smclk, smclk_en, cpu_en, dbg_en, dbg_i2c_addr_0_, dbg_i2c_addr_1_, dbg_i2c_addr_2_, dbg_i2c_addr_3_, dbg_i2c_addr_4_, dbg_i2c_addr_5_, dbg_i2c_addr_6_, dbg_i2c_broadcast_0_, dbg_i2c_broadcast_1_, dbg_i2c_broadcast_2_, dbg_i2c_broadcast_3_, dbg_i2c_broadcast_4_, dbg_i2c_broadcast_5_, dbg_i2c_broadcast_6_, dbg_i2c_scl, dbg_i2c_sda_in, dbg_uart_rxd, dco_clk, dmem_dout_0_, dmem_dout_1_, dmem_dout_2_, dmem_dout_3_, dmem_dout_4_, dmem_dout_5_, dmem_dout_6_, dmem_dout_7_, dmem_dout_8_, dmem_dout_9_, dmem_dout_10_, dmem_dout_11_, dmem_dout_12_, dmem_dout_13_, dmem_dout_14_, dmem_dout_15_, irq_0_, irq_1_, irq_2_, irq_3_, irq_4_, irq_5_, irq_6_, irq_7_, irq_8_, irq_9_, irq_10_, irq_11_, irq_12_, irq_13_, lfxt_clk, dma_addr_1_, dma_addr_2_, dma_addr_3_, dma_addr_4_, dma_addr_5_, dma_addr_6_, dma_addr_7_, dma_addr_8_, dma_addr_9_, dma_addr_10_, dma_addr_11_, dma_addr_12_, dma_addr_13_, dma_addr_14_, dma_addr_15_, dma_din_0_, dma_din_1_, dma_din_2_, dma_din_3_, dma_din_4_, dma_din_5_, dma_din_6_, dma_din_7_, dma_din_8_, dma_din_9_, dma_din_10_, dma_din_11_, dma_din_12_, dma_din_13_, dma_din_14_, dma_din_15_, dma_en, dma_priority, dma_we_0_, dma_we_1_, dma_wkup, nmi, per_dout_0_, per_dout_1_, per_dout_2_, per_dout_3_, per_dout_4_, per_dout_5_, per_dout_6_, per_dout_7_, per_dout_8_, per_dout_9_, per_dout_10_, per_dout_11_, per_dout_12_, per_dout_13_, per_dout_14_, per_dout_15_, pmem_dout_0_, pmem_dout_1_, pmem_dout_2_, pmem_dout_3_, pmem_dout_4_, pmem_dout_5_, pmem_dout_6_, pmem_dout_7_, pmem_dout_8_, pmem_dout_9_, pmem_dout_10_, pmem_dout_11_, pmem_dout_12_, pmem_dout_13_, pmem_dout_14_, pmem_dout_15_, reset_n, scan_enable, scan_mode, wkup);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire UNUSED_fe_mab_0;
  output aclk;
  output aclk_en;
  wire clock_module_0.UNUSED_cpuoff ;
  wire clock_module_0.aclk_div_0_ ;
  wire clock_module_0.aclk_div_1_ ;
  wire clock_module_0.aclk_div_2_ ;
  wire clock_module_0.bcsctl1_0_ ;
  wire clock_module_0.bcsctl1_1_ ;
  wire clock_module_0.bcsctl1_2_ ;
  wire clock_module_0.bcsctl1_3_ ;
  wire clock_module_0.bcsctl1_4_ ;
  wire clock_module_0.bcsctl1_5_ ;
  wire clock_module_0.bcsctl1_6_ ;
  wire clock_module_0.bcsctl1_7_ ;
  wire clock_module_0.bcsctl1_rd_10_ ;
  wire clock_module_0.bcsctl1_rd_11_ ;
  wire clock_module_0.bcsctl1_rd_12_ ;
  wire clock_module_0.bcsctl1_rd_13_ ;
  wire clock_module_0.bcsctl1_rd_14_ ;
  wire clock_module_0.bcsctl1_rd_15_ ;
  wire clock_module_0.bcsctl1_rd_8_ ;
  wire clock_module_0.bcsctl1_rd_9_ ;
  wire clock_module_0.bcsctl2_0_ ;
  wire clock_module_0.bcsctl2_1_ ;
  wire clock_module_0.bcsctl2_2_ ;
  wire clock_module_0.bcsctl2_3_ ;
  wire clock_module_0.bcsctl2_4_ ;
  wire clock_module_0.bcsctl2_5_ ;
  wire clock_module_0.bcsctl2_6_ ;
  wire clock_module_0.bcsctl2_7_ ;
  wire clock_module_0.bcsctl2_rd_0_ ;
  wire clock_module_0.bcsctl2_rd_1_ ;
  wire clock_module_0.bcsctl2_rd_2_ ;
  wire clock_module_0.bcsctl2_rd_3_ ;
  wire clock_module_0.bcsctl2_rd_4_ ;
  wire clock_module_0.bcsctl2_rd_5_ ;
  wire clock_module_0.bcsctl2_rd_6_ ;
  wire clock_module_0.bcsctl2_rd_7_ ;
  wire clock_module_0.dbg_cpu_reset ;
  wire clock_module_0.dbg_rst ;
  wire clock_module_0.dbg_rst_nxt ;
  wire clock_module_0.lfxt_clk_dly ;
  wire clock_module_0.lfxt_clk_s ;
  wire clock_module_0.oscoff ;
  wire clock_module_0.por ;
  wire clock_module_0.por_a ;
  wire clock_module_0.puc_a ;
  wire clock_module_0.puc_noscan_n ;
  wire clock_module_0.scg1 ;
  wire clock_module_0.smclk_div_0_ ;
  wire clock_module_0.smclk_div_1_ ;
  wire clock_module_0.smclk_div_2_ ;
  wire clock_module_0.sync_cell_lfxt_clk.data_sync_0_ ;
  wire clock_module_0.sync_cell_puc.data_in ;
  wire clock_module_0.sync_cell_puc.data_sync_0_ ;
  wire clock_module_0.sync_reset_por.data_sync_0_ ;
  wire clock_module_0.wdt_reset ;
  input cpu_en;
  wire cpu_halt_cmd;
  wire cpu_halt_st;
  wire dbg_0.UNUSED_eu_mab_0_ ;
  wire dbg_0.UNUSED_eu_mab_10_ ;
  wire dbg_0.UNUSED_eu_mab_11_ ;
  wire dbg_0.UNUSED_eu_mab_12_ ;
  wire dbg_0.UNUSED_eu_mab_13_ ;
  wire dbg_0.UNUSED_eu_mab_14_ ;
  wire dbg_0.UNUSED_eu_mab_15_ ;
  wire dbg_0.UNUSED_eu_mab_1_ ;
  wire dbg_0.UNUSED_eu_mab_2_ ;
  wire dbg_0.UNUSED_eu_mab_3_ ;
  wire dbg_0.UNUSED_eu_mab_4_ ;
  wire dbg_0.UNUSED_eu_mab_5_ ;
  wire dbg_0.UNUSED_eu_mab_6_ ;
  wire dbg_0.UNUSED_eu_mab_7_ ;
  wire dbg_0.UNUSED_eu_mab_8_ ;
  wire dbg_0.UNUSED_eu_mab_9_ ;
  wire dbg_0.UNUSED_eu_mb_en ;
  wire dbg_0.UNUSED_eu_mb_wr_0_ ;
  wire dbg_0.UNUSED_eu_mb_wr_1_ ;
  wire dbg_0.UNUSED_pc_0_ ;
  wire dbg_0.UNUSED_pc_10_ ;
  wire dbg_0.UNUSED_pc_11_ ;
  wire dbg_0.UNUSED_pc_12_ ;
  wire dbg_0.UNUSED_pc_13_ ;
  wire dbg_0.UNUSED_pc_14_ ;
  wire dbg_0.UNUSED_pc_15_ ;
  wire dbg_0.UNUSED_pc_1_ ;
  wire dbg_0.UNUSED_pc_2_ ;
  wire dbg_0.UNUSED_pc_3_ ;
  wire dbg_0.UNUSED_pc_4_ ;
  wire dbg_0.UNUSED_pc_5_ ;
  wire dbg_0.UNUSED_pc_6_ ;
  wire dbg_0.UNUSED_pc_7_ ;
  wire dbg_0.UNUSED_pc_8_ ;
  wire dbg_0.UNUSED_pc_9_ ;
  wire dbg_0.cpu_ctl_3_ ;
  wire dbg_0.cpu_ctl_4_ ;
  wire dbg_0.cpu_ctl_5_ ;
  wire dbg_0.cpu_stat_2_ ;
  wire dbg_0.cpu_stat_3_ ;
  wire dbg_0.dbg_addr_0_ ;
  wire dbg_0.dbg_addr_1_ ;
  wire dbg_0.dbg_addr_2_ ;
  wire dbg_0.dbg_addr_3_ ;
  wire dbg_0.dbg_addr_4_ ;
  wire dbg_0.dbg_addr_5_ ;
  wire dbg_0.dbg_din_0_ ;
  wire dbg_0.dbg_din_10_ ;
  wire dbg_0.dbg_din_11_ ;
  wire dbg_0.dbg_din_12_ ;
  wire dbg_0.dbg_din_13_ ;
  wire dbg_0.dbg_din_14_ ;
  wire dbg_0.dbg_din_15_ ;
  wire dbg_0.dbg_din_1_ ;
  wire dbg_0.dbg_din_2_ ;
  wire dbg_0.dbg_din_3_ ;
  wire dbg_0.dbg_din_4_ ;
  wire dbg_0.dbg_din_5_ ;
  wire dbg_0.dbg_din_6_ ;
  wire dbg_0.dbg_din_7_ ;
  wire dbg_0.dbg_din_8_ ;
  wire dbg_0.dbg_din_9_ ;
  wire dbg_0.dbg_dout_0_ ;
  wire dbg_0.dbg_dout_10_ ;
  wire dbg_0.dbg_dout_11_ ;
  wire dbg_0.dbg_dout_12_ ;
  wire dbg_0.dbg_dout_13_ ;
  wire dbg_0.dbg_dout_14_ ;
  wire dbg_0.dbg_dout_15_ ;
  wire dbg_0.dbg_dout_1_ ;
  wire dbg_0.dbg_dout_2_ ;
  wire dbg_0.dbg_dout_3_ ;
  wire dbg_0.dbg_dout_4_ ;
  wire dbg_0.dbg_dout_5_ ;
  wire dbg_0.dbg_dout_6_ ;
  wire dbg_0.dbg_dout_7_ ;
  wire dbg_0.dbg_dout_8_ ;
  wire dbg_0.dbg_dout_9_ ;
  wire dbg_0.dbg_i2c_0.dbg_bw ;
  wire dbg_0.dbg_i2c_0.dbg_rd ;
  wire dbg_0.dbg_i2c_0.dbg_state_0_ ;
  wire dbg_0.dbg_i2c_0.dbg_state_1_ ;
  wire dbg_0.dbg_i2c_0.dbg_state_2_ ;
  wire dbg_0.dbg_i2c_0.dbg_state_3_ ;
  wire dbg_0.dbg_i2c_0.dbg_state_4_ ;
  wire dbg_0.dbg_i2c_0.dbg_wr ;
  wire dbg_0.dbg_i2c_0.i2c_active_seq ;
  wire dbg_0.dbg_i2c_0.i2c_state_0_ ;
  wire dbg_0.dbg_i2c_0.i2c_state_1_ ;
  wire dbg_0.dbg_i2c_0.i2c_state_2_ ;
  wire dbg_0.dbg_i2c_0.i2c_state_3_ ;
  wire dbg_0.dbg_i2c_0.i2c_state_4_ ;
  wire dbg_0.dbg_i2c_0.i2c_state_5_ ;
  wire dbg_0.dbg_i2c_0.mem_burst ;
  wire dbg_0.dbg_i2c_0.mem_burst_end ;
  wire dbg_0.dbg_i2c_0.mem_burst_rd ;
  wire dbg_0.dbg_i2c_0.mem_burst_wr ;
  wire dbg_0.dbg_i2c_0.mem_bw ;
  wire dbg_0.dbg_i2c_0.scl ;
  wire dbg_0.dbg_i2c_0.scl_buf_0_ ;
  wire dbg_0.dbg_i2c_0.scl_buf_1_ ;
  wire dbg_0.dbg_i2c_0.scl_dly ;
  wire dbg_0.dbg_i2c_0.scl_re ;
  wire dbg_0.dbg_i2c_0.scl_re_dly_0_ ;
  wire dbg_0.dbg_i2c_0.scl_re_dly_1_ ;
  wire dbg_0.dbg_i2c_0.scl_sync ;
  wire dbg_0.dbg_i2c_0.scl_sync_n ;
  wire dbg_0.dbg_i2c_0.sda_in ;
  wire dbg_0.dbg_i2c_0.sda_in_buf_0_ ;
  wire dbg_0.dbg_i2c_0.sda_in_buf_1_ ;
  wire dbg_0.dbg_i2c_0.sda_in_dly ;
  wire dbg_0.dbg_i2c_0.sda_in_sync ;
  wire dbg_0.dbg_i2c_0.sda_in_sync_n ;
  wire dbg_0.dbg_i2c_0.shift_buf_0_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_1_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_2_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_3_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_4_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_5_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_6_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_7_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_8_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_0_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_1_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_2_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_3_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_4_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_5_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_6_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_7_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_8_ ;
  wire dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_in ;
  wire dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_sync_0_ ;
  wire dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_in ;
  wire dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_sync_0_ ;
  wire dbg_0.dbg_mem_addr_0_ ;
  wire dbg_0.dbg_mem_addr_10_ ;
  wire dbg_0.dbg_mem_addr_11_ ;
  wire dbg_0.dbg_mem_addr_12_ ;
  wire dbg_0.dbg_mem_addr_13_ ;
  wire dbg_0.dbg_mem_addr_14_ ;
  wire dbg_0.dbg_mem_addr_15_ ;
  wire dbg_0.dbg_mem_addr_1_ ;
  wire dbg_0.dbg_mem_addr_2_ ;
  wire dbg_0.dbg_mem_addr_3_ ;
  wire dbg_0.dbg_mem_addr_4_ ;
  wire dbg_0.dbg_mem_addr_5_ ;
  wire dbg_0.dbg_mem_addr_6_ ;
  wire dbg_0.dbg_mem_addr_7_ ;
  wire dbg_0.dbg_mem_addr_8_ ;
  wire dbg_0.dbg_mem_addr_9_ ;
  wire dbg_0.dbg_mem_din_0_ ;
  wire dbg_0.dbg_mem_din_10_ ;
  wire dbg_0.dbg_mem_din_11_ ;
  wire dbg_0.dbg_mem_din_12_ ;
  wire dbg_0.dbg_mem_din_13_ ;
  wire dbg_0.dbg_mem_din_14_ ;
  wire dbg_0.dbg_mem_din_15_ ;
  wire dbg_0.dbg_mem_din_1_ ;
  wire dbg_0.dbg_mem_din_2_ ;
  wire dbg_0.dbg_mem_din_3_ ;
  wire dbg_0.dbg_mem_din_4_ ;
  wire dbg_0.dbg_mem_din_5_ ;
  wire dbg_0.dbg_mem_din_6_ ;
  wire dbg_0.dbg_mem_din_7_ ;
  wire dbg_0.dbg_mem_din_8_ ;
  wire dbg_0.dbg_mem_din_9_ ;
  wire dbg_0.dbg_mem_en ;
  wire dbg_0.dbg_mem_rd ;
  wire dbg_0.dbg_mem_rd_dly ;
  wire dbg_0.dbg_mem_wr_0_ ;
  wire dbg_0.dbg_mem_wr_1_ ;
  wire dbg_0.dbg_rd_rdy ;
  wire dbg_0.dbg_reg_din_0_ ;
  wire dbg_0.dbg_reg_din_10_ ;
  wire dbg_0.dbg_reg_din_11_ ;
  wire dbg_0.dbg_reg_din_12_ ;
  wire dbg_0.dbg_reg_din_13_ ;
  wire dbg_0.dbg_reg_din_14_ ;
  wire dbg_0.dbg_reg_din_15_ ;
  wire dbg_0.dbg_reg_din_1_ ;
  wire dbg_0.dbg_reg_din_2_ ;
  wire dbg_0.dbg_reg_din_3_ ;
  wire dbg_0.dbg_reg_din_4_ ;
  wire dbg_0.dbg_reg_din_5_ ;
  wire dbg_0.dbg_reg_din_6_ ;
  wire dbg_0.dbg_reg_din_7_ ;
  wire dbg_0.dbg_reg_din_8_ ;
  wire dbg_0.dbg_reg_din_9_ ;
  wire dbg_0.dbg_reg_wr ;
  wire dbg_0.decode_noirq ;
  wire dbg_0.fe_mdb_in_0_ ;
  wire dbg_0.fe_mdb_in_10_ ;
  wire dbg_0.fe_mdb_in_11_ ;
  wire dbg_0.fe_mdb_in_12_ ;
  wire dbg_0.fe_mdb_in_13_ ;
  wire dbg_0.fe_mdb_in_14_ ;
  wire dbg_0.fe_mdb_in_15_ ;
  wire dbg_0.fe_mdb_in_1_ ;
  wire dbg_0.fe_mdb_in_2_ ;
  wire dbg_0.fe_mdb_in_3_ ;
  wire dbg_0.fe_mdb_in_4_ ;
  wire dbg_0.fe_mdb_in_5_ ;
  wire dbg_0.fe_mdb_in_6_ ;
  wire dbg_0.fe_mdb_in_7_ ;
  wire dbg_0.fe_mdb_in_8_ ;
  wire dbg_0.fe_mdb_in_9_ ;
  wire dbg_0.halt_flag ;
  wire dbg_0.inc_step_0_ ;
  wire dbg_0.inc_step_1_ ;
  wire dbg_0.istep ;
  wire dbg_0.mem_cnt_0_ ;
  wire dbg_0.mem_cnt_10_ ;
  wire dbg_0.mem_cnt_11_ ;
  wire dbg_0.mem_cnt_12_ ;
  wire dbg_0.mem_cnt_13_ ;
  wire dbg_0.mem_cnt_14_ ;
  wire dbg_0.mem_cnt_15_ ;
  wire dbg_0.mem_cnt_1_ ;
  wire dbg_0.mem_cnt_2_ ;
  wire dbg_0.mem_cnt_3_ ;
  wire dbg_0.mem_cnt_4_ ;
  wire dbg_0.mem_cnt_5_ ;
  wire dbg_0.mem_cnt_6_ ;
  wire dbg_0.mem_cnt_7_ ;
  wire dbg_0.mem_cnt_8_ ;
  wire dbg_0.mem_cnt_9_ ;
  wire dbg_0.mem_ctl_1_ ;
  wire dbg_0.mem_ctl_2_ ;
  wire dbg_0.mem_data_0_ ;
  wire dbg_0.mem_data_10_ ;
  wire dbg_0.mem_data_11_ ;
  wire dbg_0.mem_data_12_ ;
  wire dbg_0.mem_data_13_ ;
  wire dbg_0.mem_data_14_ ;
  wire dbg_0.mem_data_15_ ;
  wire dbg_0.mem_data_1_ ;
  wire dbg_0.mem_data_2_ ;
  wire dbg_0.mem_data_3_ ;
  wire dbg_0.mem_data_4_ ;
  wire dbg_0.mem_data_5_ ;
  wire dbg_0.mem_data_6_ ;
  wire dbg_0.mem_data_7_ ;
  wire dbg_0.mem_data_8_ ;
  wire dbg_0.mem_data_9_ ;
  wire dbg_0.mem_start ;
  wire dbg_0.mem_startb ;
  wire dbg_0.mem_state_0_ ;
  wire dbg_0.mem_state_1_ ;
  wire dbg_0.mem_state_2_ ;
  wire dbg_0.mem_state_3_ ;
  input dbg_en;
  output dbg_freeze;
  input dbg_i2c_addr_0_;
  input dbg_i2c_addr_1_;
  input dbg_i2c_addr_2_;
  input dbg_i2c_addr_3_;
  input dbg_i2c_addr_4_;
  input dbg_i2c_addr_5_;
  input dbg_i2c_addr_6_;
  input dbg_i2c_broadcast_0_;
  input dbg_i2c_broadcast_1_;
  input dbg_i2c_broadcast_2_;
  input dbg_i2c_broadcast_3_;
  input dbg_i2c_broadcast_4_;
  input dbg_i2c_broadcast_5_;
  input dbg_i2c_broadcast_6_;
  input dbg_i2c_scl;
  input dbg_i2c_sda_in;
  output dbg_i2c_sda_out;
  input dbg_uart_rxd;
  output dbg_uart_txd;
  input dco_clk;
  output dco_enable;
  output dco_wkup;
  input dma_addr_10_;
  input dma_addr_11_;
  input dma_addr_12_;
  input dma_addr_13_;
  input dma_addr_14_;
  input dma_addr_15_;
  input dma_addr_1_;
  input dma_addr_2_;
  input dma_addr_3_;
  input dma_addr_4_;
  input dma_addr_5_;
  input dma_addr_6_;
  input dma_addr_7_;
  input dma_addr_8_;
  input dma_addr_9_;
  input dma_din_0_;
  input dma_din_10_;
  input dma_din_11_;
  input dma_din_12_;
  input dma_din_13_;
  input dma_din_14_;
  input dma_din_15_;
  input dma_din_1_;
  input dma_din_2_;
  input dma_din_3_;
  input dma_din_4_;
  input dma_din_5_;
  input dma_din_6_;
  input dma_din_7_;
  input dma_din_8_;
  input dma_din_9_;
  output dma_dout_0_;
  output dma_dout_10_;
  output dma_dout_11_;
  output dma_dout_12_;
  output dma_dout_13_;
  output dma_dout_14_;
  output dma_dout_15_;
  output dma_dout_1_;
  output dma_dout_2_;
  output dma_dout_3_;
  output dma_dout_4_;
  output dma_dout_5_;
  output dma_dout_6_;
  output dma_dout_7_;
  output dma_dout_8_;
  output dma_dout_9_;
  input dma_en;
  input dma_priority;
  output dma_ready;
  output dma_resp;
  input dma_we_0_;
  input dma_we_1_;
  input dma_wkup;
  output dmem_addr_0_;
  output dmem_addr_10_;
  output dmem_addr_11_;
  output dmem_addr_12_;
  output dmem_addr_1_;
  output dmem_addr_2_;
  output dmem_addr_3_;
  output dmem_addr_4_;
  output dmem_addr_5_;
  output dmem_addr_6_;
  output dmem_addr_7_;
  output dmem_addr_8_;
  output dmem_addr_9_;
  output dmem_cen;
  output dmem_din_0_;
  output dmem_din_10_;
  output dmem_din_11_;
  output dmem_din_12_;
  output dmem_din_13_;
  output dmem_din_14_;
  output dmem_din_15_;
  output dmem_din_1_;
  output dmem_din_2_;
  output dmem_din_3_;
  output dmem_din_4_;
  output dmem_din_5_;
  output dmem_din_6_;
  output dmem_din_7_;
  output dmem_din_8_;
  output dmem_din_9_;
  input dmem_dout_0_;
  input dmem_dout_10_;
  input dmem_dout_11_;
  input dmem_dout_12_;
  input dmem_dout_13_;
  input dmem_dout_14_;
  input dmem_dout_15_;
  input dmem_dout_1_;
  input dmem_dout_2_;
  input dmem_dout_3_;
  input dmem_dout_4_;
  input dmem_dout_5_;
  input dmem_dout_6_;
  input dmem_dout_7_;
  input dmem_dout_8_;
  input dmem_dout_9_;
  output dmem_wen_0_;
  output dmem_wen_1_;
  wire e_state_0_;
  wire e_state_1_;
  wire e_state_2_;
  wire e_state_3_;
  wire eu_mdb_in_0_;
  wire eu_mdb_in_10_;
  wire eu_mdb_in_11_;
  wire eu_mdb_in_12_;
  wire eu_mdb_in_13_;
  wire eu_mdb_in_14_;
  wire eu_mdb_in_15_;
  wire eu_mdb_in_1_;
  wire eu_mdb_in_2_;
  wire eu_mdb_in_3_;
  wire eu_mdb_in_4_;
  wire eu_mdb_in_5_;
  wire eu_mdb_in_6_;
  wire eu_mdb_in_7_;
  wire eu_mdb_in_8_;
  wire eu_mdb_in_9_;
  wire eu_mdb_out_0_;
  wire eu_mdb_out_10_;
  wire eu_mdb_out_11_;
  wire eu_mdb_out_12_;
  wire eu_mdb_out_13_;
  wire eu_mdb_out_14_;
  wire eu_mdb_out_15_;
  wire eu_mdb_out_1_;
  wire eu_mdb_out_2_;
  wire eu_mdb_out_3_;
  wire eu_mdb_out_4_;
  wire eu_mdb_out_5_;
  wire eu_mdb_out_6_;
  wire eu_mdb_out_7_;
  wire eu_mdb_out_8_;
  wire eu_mdb_out_9_;
  wire exec_done;
  wire execution_unit_0.UNUSED_inst_ad_idx ;
  wire execution_unit_0.UNUSED_inst_ad_symb ;
  wire execution_unit_0.alu_0.N ;
  wire execution_unit_0.alu_0.UNUSED_inst_alu ;
  wire execution_unit_0.alu_0.UNUSED_inst_so_call ;
  wire execution_unit_0.alu_0.UNUSED_inst_so_push ;
  wire execution_unit_0.alu_0.UNUSED_inst_so_reti ;
  wire execution_unit_0.alu_0.Z ;
  wire execution_unit_0.alu_0.alu_out_0_ ;
  wire execution_unit_0.alu_0.alu_out_10_ ;
  wire execution_unit_0.alu_0.alu_out_11_ ;
  wire execution_unit_0.alu_0.alu_out_12_ ;
  wire execution_unit_0.alu_0.alu_out_13_ ;
  wire execution_unit_0.alu_0.alu_out_14_ ;
  wire execution_unit_0.alu_0.alu_out_15_ ;
  wire execution_unit_0.alu_0.alu_out_1_ ;
  wire execution_unit_0.alu_0.alu_out_2_ ;
  wire execution_unit_0.alu_0.alu_out_3_ ;
  wire execution_unit_0.alu_0.alu_out_4_ ;
  wire execution_unit_0.alu_0.alu_out_5_ ;
  wire execution_unit_0.alu_0.alu_out_6_ ;
  wire execution_unit_0.alu_0.alu_out_7_ ;
  wire execution_unit_0.alu_0.alu_out_8_ ;
  wire execution_unit_0.alu_0.alu_out_9_ ;
  wire execution_unit_0.alu_0.alu_shift_0_ ;
  wire execution_unit_0.alu_0.alu_shift_10_ ;
  wire execution_unit_0.alu_0.alu_shift_11_ ;
  wire execution_unit_0.alu_0.alu_shift_12_ ;
  wire execution_unit_0.alu_0.alu_shift_13_ ;
  wire execution_unit_0.alu_0.alu_shift_14_ ;
  wire execution_unit_0.alu_0.alu_shift_1_ ;
  wire execution_unit_0.alu_0.alu_shift_2_ ;
  wire execution_unit_0.alu_0.alu_shift_3_ ;
  wire execution_unit_0.alu_0.alu_shift_4_ ;
  wire execution_unit_0.alu_0.alu_shift_5_ ;
  wire execution_unit_0.alu_0.alu_shift_6_ ;
  wire execution_unit_0.alu_0.alu_shift_8_ ;
  wire execution_unit_0.alu_0.alu_shift_9_ ;
  wire execution_unit_0.alu_0.alu_stat_0_ ;
  wire execution_unit_0.alu_0.alu_stat_3_ ;
  wire execution_unit_0.alu_0.alu_stat_wr_0_ ;
  wire execution_unit_0.alu_0.alu_swpb_0_ ;
  wire execution_unit_0.alu_0.alu_swpb_8_ ;
  wire execution_unit_0.alu_0.exec_cycle ;
  wire execution_unit_0.alu_0.inst_alu_0_ ;
  wire execution_unit_0.alu_0.inst_alu_10_ ;
  wire execution_unit_0.alu_0.inst_alu_1_ ;
  wire execution_unit_0.alu_0.inst_alu_2_ ;
  wire execution_unit_0.alu_0.inst_alu_3_ ;
  wire execution_unit_0.alu_0.inst_alu_4_ ;
  wire execution_unit_0.alu_0.inst_alu_5_ ;
  wire execution_unit_0.alu_0.inst_alu_6_ ;
  wire execution_unit_0.alu_0.inst_alu_7_ ;
  wire execution_unit_0.alu_0.inst_alu_8_ ;
  wire execution_unit_0.alu_0.inst_alu_9_ ;
  wire execution_unit_0.alu_0.inst_bw ;
  wire execution_unit_0.alu_0.inst_jmp_0_ ;
  wire execution_unit_0.alu_0.inst_jmp_1_ ;
  wire execution_unit_0.alu_0.inst_jmp_2_ ;
  wire execution_unit_0.alu_0.inst_jmp_3_ ;
  wire execution_unit_0.alu_0.inst_jmp_4_ ;
  wire execution_unit_0.alu_0.inst_jmp_5_ ;
  wire execution_unit_0.alu_0.inst_jmp_6_ ;
  wire execution_unit_0.alu_0.inst_so_0_ ;
  wire execution_unit_0.alu_0.inst_so_1_ ;
  wire execution_unit_0.alu_0.inst_so_3_ ;
  wire execution_unit_0.alu_0.inst_so_7_ ;
  wire execution_unit_0.alu_0.op_dst_0_ ;
  wire execution_unit_0.alu_0.op_dst_10_ ;
  wire execution_unit_0.alu_0.op_dst_11_ ;
  wire execution_unit_0.alu_0.op_dst_12_ ;
  wire execution_unit_0.alu_0.op_dst_13_ ;
  wire execution_unit_0.alu_0.op_dst_14_ ;
  wire execution_unit_0.alu_0.op_dst_15_ ;
  wire execution_unit_0.alu_0.op_dst_1_ ;
  wire execution_unit_0.alu_0.op_dst_2_ ;
  wire execution_unit_0.alu_0.op_dst_3_ ;
  wire execution_unit_0.alu_0.op_dst_4_ ;
  wire execution_unit_0.alu_0.op_dst_5_ ;
  wire execution_unit_0.alu_0.op_dst_6_ ;
  wire execution_unit_0.alu_0.op_dst_7_ ;
  wire execution_unit_0.alu_0.op_dst_8_ ;
  wire execution_unit_0.alu_0.op_dst_9_ ;
  wire execution_unit_0.alu_0.status_0_ ;
  wire execution_unit_0.alu_0.status_1_ ;
  wire execution_unit_0.alu_0.status_2_ ;
  wire execution_unit_0.alu_0.status_3_ ;
  wire execution_unit_0.gie ;
  wire execution_unit_0.inst_ad_0_ ;
  wire execution_unit_0.inst_ad_6_ ;
  wire execution_unit_0.inst_as_0_ ;
  wire execution_unit_0.inst_as_1_ ;
  wire execution_unit_0.inst_as_2_ ;
  wire execution_unit_0.inst_as_3_ ;
  wire execution_unit_0.inst_as_4_ ;
  wire execution_unit_0.inst_as_5_ ;
  wire execution_unit_0.inst_as_6_ ;
  wire execution_unit_0.inst_as_7_ ;
  wire execution_unit_0.inst_dest_0_ ;
  wire execution_unit_0.inst_dest_10_ ;
  wire execution_unit_0.inst_dest_11_ ;
  wire execution_unit_0.inst_dest_12_ ;
  wire execution_unit_0.inst_dest_13_ ;
  wire execution_unit_0.inst_dest_14_ ;
  wire execution_unit_0.inst_dest_15_ ;
  wire execution_unit_0.inst_dest_1_ ;
  wire execution_unit_0.inst_dest_2_ ;
  wire execution_unit_0.inst_dest_3_ ;
  wire execution_unit_0.inst_dest_4_ ;
  wire execution_unit_0.inst_dest_5_ ;
  wire execution_unit_0.inst_dest_6_ ;
  wire execution_unit_0.inst_dest_7_ ;
  wire execution_unit_0.inst_dest_8_ ;
  wire execution_unit_0.inst_dest_9_ ;
  wire execution_unit_0.inst_dext_0_ ;
  wire execution_unit_0.inst_dext_10_ ;
  wire execution_unit_0.inst_dext_11_ ;
  wire execution_unit_0.inst_dext_12_ ;
  wire execution_unit_0.inst_dext_13_ ;
  wire execution_unit_0.inst_dext_14_ ;
  wire execution_unit_0.inst_dext_15_ ;
  wire execution_unit_0.inst_dext_1_ ;
  wire execution_unit_0.inst_dext_2_ ;
  wire execution_unit_0.inst_dext_3_ ;
  wire execution_unit_0.inst_dext_4_ ;
  wire execution_unit_0.inst_dext_5_ ;
  wire execution_unit_0.inst_dext_6_ ;
  wire execution_unit_0.inst_dext_7_ ;
  wire execution_unit_0.inst_dext_8_ ;
  wire execution_unit_0.inst_dext_9_ ;
  wire execution_unit_0.inst_irq_rst ;
  wire execution_unit_0.inst_mov ;
  wire execution_unit_0.inst_sext_0_ ;
  wire execution_unit_0.inst_sext_10_ ;
  wire execution_unit_0.inst_sext_11_ ;
  wire execution_unit_0.inst_sext_12_ ;
  wire execution_unit_0.inst_sext_13_ ;
  wire execution_unit_0.inst_sext_14_ ;
  wire execution_unit_0.inst_sext_15_ ;
  wire execution_unit_0.inst_sext_1_ ;
  wire execution_unit_0.inst_sext_2_ ;
  wire execution_unit_0.inst_sext_3_ ;
  wire execution_unit_0.inst_sext_4_ ;
  wire execution_unit_0.inst_sext_5_ ;
  wire execution_unit_0.inst_sext_6_ ;
  wire execution_unit_0.inst_sext_7_ ;
  wire execution_unit_0.inst_sext_8_ ;
  wire execution_unit_0.inst_sext_9_ ;
  wire execution_unit_0.inst_src_0_ ;
  wire execution_unit_0.inst_src_10_ ;
  wire execution_unit_0.inst_src_11_ ;
  wire execution_unit_0.inst_src_12_ ;
  wire execution_unit_0.inst_src_13_ ;
  wire execution_unit_0.inst_src_14_ ;
  wire execution_unit_0.inst_src_15_ ;
  wire execution_unit_0.inst_src_1_ ;
  wire execution_unit_0.inst_src_2_ ;
  wire execution_unit_0.inst_src_3_ ;
  wire execution_unit_0.inst_src_4_ ;
  wire execution_unit_0.inst_src_5_ ;
  wire execution_unit_0.inst_src_6_ ;
  wire execution_unit_0.inst_src_7_ ;
  wire execution_unit_0.inst_src_8_ ;
  wire execution_unit_0.inst_src_9_ ;
  wire execution_unit_0.inst_type_0_ ;
  wire execution_unit_0.inst_type_1_ ;
  wire execution_unit_0.inst_type_2_ ;
  wire execution_unit_0.mab_lsb ;
  wire execution_unit_0.mdb_in_buf_0_ ;
  wire execution_unit_0.mdb_in_buf_10_ ;
  wire execution_unit_0.mdb_in_buf_11_ ;
  wire execution_unit_0.mdb_in_buf_12_ ;
  wire execution_unit_0.mdb_in_buf_13_ ;
  wire execution_unit_0.mdb_in_buf_14_ ;
  wire execution_unit_0.mdb_in_buf_15_ ;
  wire execution_unit_0.mdb_in_buf_1_ ;
  wire execution_unit_0.mdb_in_buf_2_ ;
  wire execution_unit_0.mdb_in_buf_3_ ;
  wire execution_unit_0.mdb_in_buf_4_ ;
  wire execution_unit_0.mdb_in_buf_5_ ;
  wire execution_unit_0.mdb_in_buf_6_ ;
  wire execution_unit_0.mdb_in_buf_7_ ;
  wire execution_unit_0.mdb_in_buf_8_ ;
  wire execution_unit_0.mdb_in_buf_9_ ;
  wire execution_unit_0.mdb_in_buf_en ;
  wire execution_unit_0.mdb_in_buf_valid ;
  wire execution_unit_0.mdb_out_nxt_10_ ;
  wire execution_unit_0.mdb_out_nxt_11_ ;
  wire execution_unit_0.mdb_out_nxt_12_ ;
  wire execution_unit_0.mdb_out_nxt_13_ ;
  wire execution_unit_0.mdb_out_nxt_14_ ;
  wire execution_unit_0.mdb_out_nxt_15_ ;
  wire execution_unit_0.mdb_out_nxt_8_ ;
  wire execution_unit_0.mdb_out_nxt_9_ ;
  wire execution_unit_0.pc_nxt_10_ ;
  wire execution_unit_0.pc_nxt_11_ ;
  wire execution_unit_0.pc_nxt_12_ ;
  wire execution_unit_0.pc_nxt_13_ ;
  wire execution_unit_0.pc_nxt_14_ ;
  wire execution_unit_0.pc_nxt_15_ ;
  wire execution_unit_0.pc_nxt_1_ ;
  wire execution_unit_0.pc_nxt_2_ ;
  wire execution_unit_0.pc_nxt_3_ ;
  wire execution_unit_0.pc_nxt_4_ ;
  wire execution_unit_0.pc_nxt_5_ ;
  wire execution_unit_0.pc_nxt_6_ ;
  wire execution_unit_0.pc_nxt_7_ ;
  wire execution_unit_0.pc_nxt_8_ ;
  wire execution_unit_0.pc_nxt_9_ ;
  wire execution_unit_0.pc_sw_10_ ;
  wire execution_unit_0.pc_sw_11_ ;
  wire execution_unit_0.pc_sw_12_ ;
  wire execution_unit_0.pc_sw_13_ ;
  wire execution_unit_0.pc_sw_14_ ;
  wire execution_unit_0.pc_sw_15_ ;
  wire execution_unit_0.pc_sw_8_ ;
  wire execution_unit_0.pc_sw_9_ ;
  wire execution_unit_0.pc_sw_wr ;
  wire execution_unit_0.reg_dest_wr ;
  wire execution_unit_0.reg_incr ;
  wire execution_unit_0.reg_pc_call ;
  wire execution_unit_0.reg_sp_wr ;
  wire execution_unit_0.reg_sr_clr ;
  wire execution_unit_0.reg_sr_wr ;
  wire execution_unit_0.reg_src_0_ ;
  wire execution_unit_0.reg_src_10_ ;
  wire execution_unit_0.reg_src_11_ ;
  wire execution_unit_0.reg_src_12_ ;
  wire execution_unit_0.reg_src_13_ ;
  wire execution_unit_0.reg_src_14_ ;
  wire execution_unit_0.reg_src_15_ ;
  wire execution_unit_0.reg_src_1_ ;
  wire execution_unit_0.reg_src_2_ ;
  wire execution_unit_0.reg_src_3_ ;
  wire execution_unit_0.reg_src_4_ ;
  wire execution_unit_0.reg_src_5_ ;
  wire execution_unit_0.reg_src_6_ ;
  wire execution_unit_0.reg_src_7_ ;
  wire execution_unit_0.reg_src_8_ ;
  wire execution_unit_0.reg_src_9_ ;
  wire execution_unit_0.register_file_0.r10_0_ ;
  wire execution_unit_0.register_file_0.r10_10_ ;
  wire execution_unit_0.register_file_0.r10_11_ ;
  wire execution_unit_0.register_file_0.r10_12_ ;
  wire execution_unit_0.register_file_0.r10_13_ ;
  wire execution_unit_0.register_file_0.r10_14_ ;
  wire execution_unit_0.register_file_0.r10_15_ ;
  wire execution_unit_0.register_file_0.r10_1_ ;
  wire execution_unit_0.register_file_0.r10_2_ ;
  wire execution_unit_0.register_file_0.r10_3_ ;
  wire execution_unit_0.register_file_0.r10_4_ ;
  wire execution_unit_0.register_file_0.r10_5_ ;
  wire execution_unit_0.register_file_0.r10_6_ ;
  wire execution_unit_0.register_file_0.r10_7_ ;
  wire execution_unit_0.register_file_0.r10_8_ ;
  wire execution_unit_0.register_file_0.r10_9_ ;
  wire execution_unit_0.register_file_0.r11_0_ ;
  wire execution_unit_0.register_file_0.r11_10_ ;
  wire execution_unit_0.register_file_0.r11_11_ ;
  wire execution_unit_0.register_file_0.r11_12_ ;
  wire execution_unit_0.register_file_0.r11_13_ ;
  wire execution_unit_0.register_file_0.r11_14_ ;
  wire execution_unit_0.register_file_0.r11_15_ ;
  wire execution_unit_0.register_file_0.r11_1_ ;
  wire execution_unit_0.register_file_0.r11_2_ ;
  wire execution_unit_0.register_file_0.r11_3_ ;
  wire execution_unit_0.register_file_0.r11_4_ ;
  wire execution_unit_0.register_file_0.r11_5_ ;
  wire execution_unit_0.register_file_0.r11_6_ ;
  wire execution_unit_0.register_file_0.r11_7_ ;
  wire execution_unit_0.register_file_0.r11_8_ ;
  wire execution_unit_0.register_file_0.r11_9_ ;
  wire execution_unit_0.register_file_0.r12_0_ ;
  wire execution_unit_0.register_file_0.r12_10_ ;
  wire execution_unit_0.register_file_0.r12_11_ ;
  wire execution_unit_0.register_file_0.r12_12_ ;
  wire execution_unit_0.register_file_0.r12_13_ ;
  wire execution_unit_0.register_file_0.r12_14_ ;
  wire execution_unit_0.register_file_0.r12_15_ ;
  wire execution_unit_0.register_file_0.r12_1_ ;
  wire execution_unit_0.register_file_0.r12_2_ ;
  wire execution_unit_0.register_file_0.r12_3_ ;
  wire execution_unit_0.register_file_0.r12_4_ ;
  wire execution_unit_0.register_file_0.r12_5_ ;
  wire execution_unit_0.register_file_0.r12_6_ ;
  wire execution_unit_0.register_file_0.r12_7_ ;
  wire execution_unit_0.register_file_0.r12_8_ ;
  wire execution_unit_0.register_file_0.r12_9_ ;
  wire execution_unit_0.register_file_0.r13_0_ ;
  wire execution_unit_0.register_file_0.r13_10_ ;
  wire execution_unit_0.register_file_0.r13_11_ ;
  wire execution_unit_0.register_file_0.r13_12_ ;
  wire execution_unit_0.register_file_0.r13_13_ ;
  wire execution_unit_0.register_file_0.r13_14_ ;
  wire execution_unit_0.register_file_0.r13_15_ ;
  wire execution_unit_0.register_file_0.r13_1_ ;
  wire execution_unit_0.register_file_0.r13_2_ ;
  wire execution_unit_0.register_file_0.r13_3_ ;
  wire execution_unit_0.register_file_0.r13_4_ ;
  wire execution_unit_0.register_file_0.r13_5_ ;
  wire execution_unit_0.register_file_0.r13_6_ ;
  wire execution_unit_0.register_file_0.r13_7_ ;
  wire execution_unit_0.register_file_0.r13_8_ ;
  wire execution_unit_0.register_file_0.r13_9_ ;
  wire execution_unit_0.register_file_0.r14_0_ ;
  wire execution_unit_0.register_file_0.r14_10_ ;
  wire execution_unit_0.register_file_0.r14_11_ ;
  wire execution_unit_0.register_file_0.r14_12_ ;
  wire execution_unit_0.register_file_0.r14_13_ ;
  wire execution_unit_0.register_file_0.r14_14_ ;
  wire execution_unit_0.register_file_0.r14_15_ ;
  wire execution_unit_0.register_file_0.r14_1_ ;
  wire execution_unit_0.register_file_0.r14_2_ ;
  wire execution_unit_0.register_file_0.r14_3_ ;
  wire execution_unit_0.register_file_0.r14_4_ ;
  wire execution_unit_0.register_file_0.r14_5_ ;
  wire execution_unit_0.register_file_0.r14_6_ ;
  wire execution_unit_0.register_file_0.r14_7_ ;
  wire execution_unit_0.register_file_0.r14_8_ ;
  wire execution_unit_0.register_file_0.r14_9_ ;
  wire execution_unit_0.register_file_0.r15_0_ ;
  wire execution_unit_0.register_file_0.r15_10_ ;
  wire execution_unit_0.register_file_0.r15_11_ ;
  wire execution_unit_0.register_file_0.r15_12_ ;
  wire execution_unit_0.register_file_0.r15_13_ ;
  wire execution_unit_0.register_file_0.r15_14_ ;
  wire execution_unit_0.register_file_0.r15_15_ ;
  wire execution_unit_0.register_file_0.r15_1_ ;
  wire execution_unit_0.register_file_0.r15_2_ ;
  wire execution_unit_0.register_file_0.r15_3_ ;
  wire execution_unit_0.register_file_0.r15_4_ ;
  wire execution_unit_0.register_file_0.r15_5_ ;
  wire execution_unit_0.register_file_0.r15_6_ ;
  wire execution_unit_0.register_file_0.r15_7_ ;
  wire execution_unit_0.register_file_0.r15_8_ ;
  wire execution_unit_0.register_file_0.r15_9_ ;
  wire execution_unit_0.register_file_0.r1_0_ ;
  wire execution_unit_0.register_file_0.r1_10_ ;
  wire execution_unit_0.register_file_0.r1_11_ ;
  wire execution_unit_0.register_file_0.r1_12_ ;
  wire execution_unit_0.register_file_0.r1_13_ ;
  wire execution_unit_0.register_file_0.r1_14_ ;
  wire execution_unit_0.register_file_0.r1_15_ ;
  wire execution_unit_0.register_file_0.r1_1_ ;
  wire execution_unit_0.register_file_0.r1_2_ ;
  wire execution_unit_0.register_file_0.r1_3_ ;
  wire execution_unit_0.register_file_0.r1_4_ ;
  wire execution_unit_0.register_file_0.r1_5_ ;
  wire execution_unit_0.register_file_0.r1_6_ ;
  wire execution_unit_0.register_file_0.r1_7_ ;
  wire execution_unit_0.register_file_0.r1_8_ ;
  wire execution_unit_0.register_file_0.r1_9_ ;
  wire execution_unit_0.register_file_0.r2_4_ ;
  wire execution_unit_0.register_file_0.r3_0_ ;
  wire execution_unit_0.register_file_0.r3_10_ ;
  wire execution_unit_0.register_file_0.r3_11_ ;
  wire execution_unit_0.register_file_0.r3_12_ ;
  wire execution_unit_0.register_file_0.r3_13_ ;
  wire execution_unit_0.register_file_0.r3_14_ ;
  wire execution_unit_0.register_file_0.r3_15_ ;
  wire execution_unit_0.register_file_0.r3_1_ ;
  wire execution_unit_0.register_file_0.r3_2_ ;
  wire execution_unit_0.register_file_0.r3_3_ ;
  wire execution_unit_0.register_file_0.r3_4_ ;
  wire execution_unit_0.register_file_0.r3_5_ ;
  wire execution_unit_0.register_file_0.r3_6_ ;
  wire execution_unit_0.register_file_0.r3_7_ ;
  wire execution_unit_0.register_file_0.r3_8_ ;
  wire execution_unit_0.register_file_0.r3_9_ ;
  wire execution_unit_0.register_file_0.r4_0_ ;
  wire execution_unit_0.register_file_0.r4_10_ ;
  wire execution_unit_0.register_file_0.r4_11_ ;
  wire execution_unit_0.register_file_0.r4_12_ ;
  wire execution_unit_0.register_file_0.r4_13_ ;
  wire execution_unit_0.register_file_0.r4_14_ ;
  wire execution_unit_0.register_file_0.r4_15_ ;
  wire execution_unit_0.register_file_0.r4_1_ ;
  wire execution_unit_0.register_file_0.r4_2_ ;
  wire execution_unit_0.register_file_0.r4_3_ ;
  wire execution_unit_0.register_file_0.r4_4_ ;
  wire execution_unit_0.register_file_0.r4_5_ ;
  wire execution_unit_0.register_file_0.r4_6_ ;
  wire execution_unit_0.register_file_0.r4_7_ ;
  wire execution_unit_0.register_file_0.r4_8_ ;
  wire execution_unit_0.register_file_0.r4_9_ ;
  wire execution_unit_0.register_file_0.r5_0_ ;
  wire execution_unit_0.register_file_0.r5_10_ ;
  wire execution_unit_0.register_file_0.r5_11_ ;
  wire execution_unit_0.register_file_0.r5_12_ ;
  wire execution_unit_0.register_file_0.r5_13_ ;
  wire execution_unit_0.register_file_0.r5_14_ ;
  wire execution_unit_0.register_file_0.r5_15_ ;
  wire execution_unit_0.register_file_0.r5_1_ ;
  wire execution_unit_0.register_file_0.r5_2_ ;
  wire execution_unit_0.register_file_0.r5_3_ ;
  wire execution_unit_0.register_file_0.r5_4_ ;
  wire execution_unit_0.register_file_0.r5_5_ ;
  wire execution_unit_0.register_file_0.r5_6_ ;
  wire execution_unit_0.register_file_0.r5_7_ ;
  wire execution_unit_0.register_file_0.r5_8_ ;
  wire execution_unit_0.register_file_0.r5_9_ ;
  wire execution_unit_0.register_file_0.r6_0_ ;
  wire execution_unit_0.register_file_0.r6_10_ ;
  wire execution_unit_0.register_file_0.r6_11_ ;
  wire execution_unit_0.register_file_0.r6_12_ ;
  wire execution_unit_0.register_file_0.r6_13_ ;
  wire execution_unit_0.register_file_0.r6_14_ ;
  wire execution_unit_0.register_file_0.r6_15_ ;
  wire execution_unit_0.register_file_0.r6_1_ ;
  wire execution_unit_0.register_file_0.r6_2_ ;
  wire execution_unit_0.register_file_0.r6_3_ ;
  wire execution_unit_0.register_file_0.r6_4_ ;
  wire execution_unit_0.register_file_0.r6_5_ ;
  wire execution_unit_0.register_file_0.r6_6_ ;
  wire execution_unit_0.register_file_0.r6_7_ ;
  wire execution_unit_0.register_file_0.r6_8_ ;
  wire execution_unit_0.register_file_0.r6_9_ ;
  wire execution_unit_0.register_file_0.r7_0_ ;
  wire execution_unit_0.register_file_0.r7_10_ ;
  wire execution_unit_0.register_file_0.r7_11_ ;
  wire execution_unit_0.register_file_0.r7_12_ ;
  wire execution_unit_0.register_file_0.r7_13_ ;
  wire execution_unit_0.register_file_0.r7_14_ ;
  wire execution_unit_0.register_file_0.r7_15_ ;
  wire execution_unit_0.register_file_0.r7_1_ ;
  wire execution_unit_0.register_file_0.r7_2_ ;
  wire execution_unit_0.register_file_0.r7_3_ ;
  wire execution_unit_0.register_file_0.r7_4_ ;
  wire execution_unit_0.register_file_0.r7_5_ ;
  wire execution_unit_0.register_file_0.r7_6_ ;
  wire execution_unit_0.register_file_0.r7_7_ ;
  wire execution_unit_0.register_file_0.r7_8_ ;
  wire execution_unit_0.register_file_0.r7_9_ ;
  wire execution_unit_0.register_file_0.r8_0_ ;
  wire execution_unit_0.register_file_0.r8_10_ ;
  wire execution_unit_0.register_file_0.r8_11_ ;
  wire execution_unit_0.register_file_0.r8_12_ ;
  wire execution_unit_0.register_file_0.r8_13_ ;
  wire execution_unit_0.register_file_0.r8_14_ ;
  wire execution_unit_0.register_file_0.r8_15_ ;
  wire execution_unit_0.register_file_0.r8_1_ ;
  wire execution_unit_0.register_file_0.r8_2_ ;
  wire execution_unit_0.register_file_0.r8_3_ ;
  wire execution_unit_0.register_file_0.r8_4_ ;
  wire execution_unit_0.register_file_0.r8_5_ ;
  wire execution_unit_0.register_file_0.r8_6_ ;
  wire execution_unit_0.register_file_0.r8_7_ ;
  wire execution_unit_0.register_file_0.r8_8_ ;
  wire execution_unit_0.register_file_0.r8_9_ ;
  wire execution_unit_0.register_file_0.r9_0_ ;
  wire execution_unit_0.register_file_0.r9_10_ ;
  wire execution_unit_0.register_file_0.r9_11_ ;
  wire execution_unit_0.register_file_0.r9_12_ ;
  wire execution_unit_0.register_file_0.r9_13_ ;
  wire execution_unit_0.register_file_0.r9_14_ ;
  wire execution_unit_0.register_file_0.r9_15_ ;
  wire execution_unit_0.register_file_0.r9_1_ ;
  wire execution_unit_0.register_file_0.r9_2_ ;
  wire execution_unit_0.register_file_0.r9_3_ ;
  wire execution_unit_0.register_file_0.r9_4_ ;
  wire execution_unit_0.register_file_0.r9_5_ ;
  wire execution_unit_0.register_file_0.r9_6_ ;
  wire execution_unit_0.register_file_0.r9_7_ ;
  wire execution_unit_0.register_file_0.r9_8_ ;
  wire execution_unit_0.register_file_0.r9_9_ ;
  wire fe_mb_en;
  wire fe_pmem_wait;
  wire frontend_0.e_state_nxt_0_ ;
  wire frontend_0.e_state_nxt_1_ ;
  wire frontend_0.e_state_nxt_2_ ;
  wire frontend_0.e_state_nxt_3_ ;
  wire frontend_0.exec_dext_rdy ;
  wire frontend_0.exec_dst_wr ;
  wire frontend_0.exec_jmp ;
  wire frontend_0.exec_src_wr ;
  wire frontend_0.i_state_0_ ;
  wire frontend_0.i_state_1_ ;
  wire frontend_0.i_state_2_ ;
  wire frontend_0.i_state_3_ ;
  wire frontend_0.i_state_4_ ;
  wire frontend_0.i_state_5_ ;
  wire frontend_0.inst_dest_bin_0_ ;
  wire frontend_0.inst_dest_bin_1_ ;
  wire frontend_0.inst_dest_bin_2_ ;
  wire frontend_0.inst_dest_bin_3_ ;
  wire frontend_0.inst_jmp_bin_0_ ;
  wire frontend_0.inst_jmp_bin_1_ ;
  wire frontend_0.inst_jmp_bin_2_ ;
  wire frontend_0.inst_src_bin_0_ ;
  wire frontend_0.inst_src_bin_1_ ;
  wire frontend_0.inst_src_bin_2_ ;
  wire frontend_0.inst_src_bin_3_ ;
  wire frontend_0.inst_sz_0_ ;
  wire frontend_0.inst_sz_1_ ;
  wire frontend_0.irq_addr_1_ ;
  wire frontend_0.irq_addr_2_ ;
  wire frontend_0.irq_addr_3_ ;
  wire frontend_0.irq_addr_4_ ;
  wire frontend_0.irq_addr_5_ ;
  wire frontend_0.irq_addr_6_ ;
  wire frontend_0.pmem_busy ;
  wire frontend_0.wdt_irq ;
  input irq_0_;
  input irq_10_;
  input irq_11_;
  input irq_12_;
  input irq_13_;
  input irq_1_;
  input irq_2_;
  input irq_3_;
  input irq_4_;
  input irq_5_;
  input irq_6_;
  input irq_7_;
  input irq_8_;
  input irq_9_;
  output irq_acc_0_;
  output irq_acc_10_;
  output irq_acc_11_;
  output irq_acc_12_;
  output irq_acc_13_;
  output irq_acc_1_;
  output irq_acc_2_;
  output irq_acc_3_;
  output irq_acc_4_;
  output irq_acc_5_;
  output irq_acc_6_;
  output irq_acc_7_;
  output irq_acc_8_;
  output irq_acc_9_;
  input lfxt_clk;
  output lfxt_enable;
  output lfxt_wkup;
  output mclk;
  wire mem_backbone_0.eu_mdb_in_sel_0_ ;
  wire mem_backbone_0.eu_mdb_in_sel_1_ ;
  wire mem_backbone_0.eu_per_en ;
  wire mem_backbone_0.eu_pmem_en ;
  wire mem_backbone_0.ext_mem_din_sel_0_ ;
  wire mem_backbone_0.ext_mem_din_sel_1_ ;
  wire mem_backbone_0.ext_per_en ;
  wire mem_backbone_0.ext_pmem_en ;
  wire mem_backbone_0.fe_pmem_en ;
  wire mem_backbone_0.fe_pmem_en_dly ;
  wire mem_backbone_0.per_dout_0_ ;
  wire mem_backbone_0.per_dout_10_ ;
  wire mem_backbone_0.per_dout_11_ ;
  wire mem_backbone_0.per_dout_12_ ;
  wire mem_backbone_0.per_dout_13_ ;
  wire mem_backbone_0.per_dout_14_ ;
  wire mem_backbone_0.per_dout_15_ ;
  wire mem_backbone_0.per_dout_1_ ;
  wire mem_backbone_0.per_dout_2_ ;
  wire mem_backbone_0.per_dout_3_ ;
  wire mem_backbone_0.per_dout_4_ ;
  wire mem_backbone_0.per_dout_5_ ;
  wire mem_backbone_0.per_dout_6_ ;
  wire mem_backbone_0.per_dout_7_ ;
  wire mem_backbone_0.per_dout_8_ ;
  wire mem_backbone_0.per_dout_9_ ;
  wire mem_backbone_0.per_dout_val_0_ ;
  wire mem_backbone_0.per_dout_val_10_ ;
  wire mem_backbone_0.per_dout_val_11_ ;
  wire mem_backbone_0.per_dout_val_12_ ;
  wire mem_backbone_0.per_dout_val_13_ ;
  wire mem_backbone_0.per_dout_val_14_ ;
  wire mem_backbone_0.per_dout_val_15_ ;
  wire mem_backbone_0.per_dout_val_1_ ;
  wire mem_backbone_0.per_dout_val_2_ ;
  wire mem_backbone_0.per_dout_val_3_ ;
  wire mem_backbone_0.per_dout_val_4_ ;
  wire mem_backbone_0.per_dout_val_5_ ;
  wire mem_backbone_0.per_dout_val_6_ ;
  wire mem_backbone_0.per_dout_val_7_ ;
  wire mem_backbone_0.per_dout_val_8_ ;
  wire mem_backbone_0.per_dout_val_9_ ;
  wire mem_backbone_0.pmem_dout_bckup_0_ ;
  wire mem_backbone_0.pmem_dout_bckup_10_ ;
  wire mem_backbone_0.pmem_dout_bckup_11_ ;
  wire mem_backbone_0.pmem_dout_bckup_12_ ;
  wire mem_backbone_0.pmem_dout_bckup_13_ ;
  wire mem_backbone_0.pmem_dout_bckup_14_ ;
  wire mem_backbone_0.pmem_dout_bckup_15_ ;
  wire mem_backbone_0.pmem_dout_bckup_1_ ;
  wire mem_backbone_0.pmem_dout_bckup_2_ ;
  wire mem_backbone_0.pmem_dout_bckup_3_ ;
  wire mem_backbone_0.pmem_dout_bckup_4_ ;
  wire mem_backbone_0.pmem_dout_bckup_5_ ;
  wire mem_backbone_0.pmem_dout_bckup_6_ ;
  wire mem_backbone_0.pmem_dout_bckup_7_ ;
  wire mem_backbone_0.pmem_dout_bckup_8_ ;
  wire mem_backbone_0.pmem_dout_bckup_9_ ;
  wire mem_backbone_0.pmem_dout_bckup_sel ;
  wire multiplier_0.acc_sel ;
  wire multiplier_0.cycle_0_ ;
  wire multiplier_0.cycle_1_ ;
  wire multiplier_0.op1_0_ ;
  wire multiplier_0.op1_10_ ;
  wire multiplier_0.op1_11_ ;
  wire multiplier_0.op1_12_ ;
  wire multiplier_0.op1_13_ ;
  wire multiplier_0.op1_14_ ;
  wire multiplier_0.op1_15_ ;
  wire multiplier_0.op1_1_ ;
  wire multiplier_0.op1_2_ ;
  wire multiplier_0.op1_3_ ;
  wire multiplier_0.op1_4_ ;
  wire multiplier_0.op1_5_ ;
  wire multiplier_0.op1_6_ ;
  wire multiplier_0.op1_7_ ;
  wire multiplier_0.op1_8_ ;
  wire multiplier_0.op1_9_ ;
  wire multiplier_0.op2_0_ ;
  wire multiplier_0.op2_10_ ;
  wire multiplier_0.op2_11_ ;
  wire multiplier_0.op2_12_ ;
  wire multiplier_0.op2_13_ ;
  wire multiplier_0.op2_14_ ;
  wire multiplier_0.op2_15_ ;
  wire multiplier_0.op2_1_ ;
  wire multiplier_0.op2_2_ ;
  wire multiplier_0.op2_3_ ;
  wire multiplier_0.op2_4_ ;
  wire multiplier_0.op2_5_ ;
  wire multiplier_0.op2_6_ ;
  wire multiplier_0.op2_7_ ;
  wire multiplier_0.op2_8_ ;
  wire multiplier_0.op2_9_ ;
  wire multiplier_0.op2_wr ;
  wire multiplier_0.per_dout_0_ ;
  wire multiplier_0.per_dout_10_ ;
  wire multiplier_0.per_dout_11_ ;
  wire multiplier_0.per_dout_12_ ;
  wire multiplier_0.per_dout_13_ ;
  wire multiplier_0.per_dout_14_ ;
  wire multiplier_0.per_dout_15_ ;
  wire multiplier_0.per_dout_1_ ;
  wire multiplier_0.per_dout_2_ ;
  wire multiplier_0.per_dout_3_ ;
  wire multiplier_0.per_dout_4_ ;
  wire multiplier_0.per_dout_5_ ;
  wire multiplier_0.per_dout_6_ ;
  wire multiplier_0.per_dout_7_ ;
  wire multiplier_0.per_dout_8_ ;
  wire multiplier_0.per_dout_9_ ;
  wire multiplier_0.reshi_0_ ;
  wire multiplier_0.reshi_10_ ;
  wire multiplier_0.reshi_11_ ;
  wire multiplier_0.reshi_12_ ;
  wire multiplier_0.reshi_13_ ;
  wire multiplier_0.reshi_14_ ;
  wire multiplier_0.reshi_15_ ;
  wire multiplier_0.reshi_1_ ;
  wire multiplier_0.reshi_2_ ;
  wire multiplier_0.reshi_3_ ;
  wire multiplier_0.reshi_4_ ;
  wire multiplier_0.reshi_5_ ;
  wire multiplier_0.reshi_6_ ;
  wire multiplier_0.reshi_7_ ;
  wire multiplier_0.reshi_8_ ;
  wire multiplier_0.reshi_9_ ;
  wire multiplier_0.reslo_0_ ;
  wire multiplier_0.reslo_10_ ;
  wire multiplier_0.reslo_11_ ;
  wire multiplier_0.reslo_12_ ;
  wire multiplier_0.reslo_13_ ;
  wire multiplier_0.reslo_14_ ;
  wire multiplier_0.reslo_15_ ;
  wire multiplier_0.reslo_1_ ;
  wire multiplier_0.reslo_2_ ;
  wire multiplier_0.reslo_3_ ;
  wire multiplier_0.reslo_4_ ;
  wire multiplier_0.reslo_5_ ;
  wire multiplier_0.reslo_6_ ;
  wire multiplier_0.reslo_7_ ;
  wire multiplier_0.reslo_8_ ;
  wire multiplier_0.reslo_9_ ;
  wire multiplier_0.sign_sel ;
  wire multiplier_0.sumext_0_ ;
  wire multiplier_0.sumext_10_ ;
  input nmi;
  output per_addr_0_;
  output per_addr_10_;
  output per_addr_11_;
  output per_addr_12_;
  output per_addr_13_;
  output per_addr_1_;
  output per_addr_2_;
  output per_addr_3_;
  output per_addr_4_;
  output per_addr_5_;
  output per_addr_6_;
  output per_addr_7_;
  output per_addr_8_;
  output per_addr_9_;
  output per_din_0_;
  output per_din_10_;
  output per_din_11_;
  output per_din_12_;
  output per_din_13_;
  output per_din_14_;
  output per_din_15_;
  output per_din_1_;
  output per_din_2_;
  output per_din_3_;
  output per_din_4_;
  output per_din_5_;
  output per_din_6_;
  output per_din_7_;
  output per_din_8_;
  output per_din_9_;
  input per_dout_0_;
  input per_dout_10_;
  input per_dout_11_;
  input per_dout_12_;
  input per_dout_13_;
  input per_dout_14_;
  input per_dout_15_;
  input per_dout_1_;
  input per_dout_2_;
  input per_dout_3_;
  input per_dout_4_;
  input per_dout_5_;
  input per_dout_6_;
  input per_dout_7_;
  input per_dout_8_;
  input per_dout_9_;
  wire per_dout_sfr_0_;
  wire per_dout_sfr_10_;
  wire per_dout_sfr_11_;
  wire per_dout_sfr_12_;
  wire per_dout_sfr_13_;
  wire per_dout_sfr_14_;
  wire per_dout_sfr_15_;
  wire per_dout_sfr_1_;
  wire per_dout_sfr_2_;
  wire per_dout_sfr_3_;
  wire per_dout_sfr_4_;
  wire per_dout_sfr_5_;
  wire per_dout_sfr_6_;
  wire per_dout_sfr_7_;
  wire per_dout_sfr_8_;
  wire per_dout_sfr_9_;
  wire per_dout_wdog_0_;
  wire per_dout_wdog_11_;
  wire per_dout_wdog_1_;
  wire per_dout_wdog_2_;
  wire per_dout_wdog_3_;
  wire per_dout_wdog_4_;
  wire per_dout_wdog_5_;
  wire per_dout_wdog_6_;
  wire per_dout_wdog_7_;
  output per_en;
  output per_we_0_;
  output per_we_1_;
  output pmem_addr_0_;
  output pmem_addr_10_;
  output pmem_addr_11_;
  output pmem_addr_12_;
  output pmem_addr_13_;
  output pmem_addr_1_;
  output pmem_addr_2_;
  output pmem_addr_3_;
  output pmem_addr_4_;
  output pmem_addr_5_;
  output pmem_addr_6_;
  output pmem_addr_7_;
  output pmem_addr_8_;
  output pmem_addr_9_;
  output pmem_cen;
  output pmem_din_0_;
  output pmem_din_10_;
  output pmem_din_11_;
  output pmem_din_12_;
  output pmem_din_13_;
  output pmem_din_14_;
  output pmem_din_15_;
  output pmem_din_1_;
  output pmem_din_2_;
  output pmem_din_3_;
  output pmem_din_4_;
  output pmem_din_5_;
  output pmem_din_6_;
  output pmem_din_7_;
  output pmem_din_8_;
  output pmem_din_9_;
  input pmem_dout_0_;
  input pmem_dout_10_;
  input pmem_dout_11_;
  input pmem_dout_12_;
  input pmem_dout_13_;
  input pmem_dout_14_;
  input pmem_dout_15_;
  input pmem_dout_1_;
  input pmem_dout_2_;
  input pmem_dout_3_;
  input pmem_dout_4_;
  input pmem_dout_5_;
  input pmem_dout_6_;
  input pmem_dout_7_;
  input pmem_dout_8_;
  input pmem_dout_9_;
  output pmem_wen_0_;
  output pmem_wen_1_;
  output puc_rst;
  input reset_n;
  input scan_enable;
  input scan_mode;
  wire sfr_0.UNUSED_wdtnmies ;
  wire sfr_0.ie1_0_ ;
  wire sfr_0.ifg1_0_ ;
  wire sfr_0.wdtifg_sw_clr ;
  wire sfr_0.wdtifg_sw_set ;
  output smclk;
  output smclk_en;
  wire watchdog_0.wdtcnt_0_ ;
  wire watchdog_0.wdtcnt_10_ ;
  wire watchdog_0.wdtcnt_11_ ;
  wire watchdog_0.wdtcnt_12_ ;
  wire watchdog_0.wdtcnt_13_ ;
  wire watchdog_0.wdtcnt_14_ ;
  wire watchdog_0.wdtcnt_15_ ;
  wire watchdog_0.wdtcnt_1_ ;
  wire watchdog_0.wdtcnt_2_ ;
  wire watchdog_0.wdtcnt_3_ ;
  wire watchdog_0.wdtcnt_4_ ;
  wire watchdog_0.wdtcnt_5_ ;
  wire watchdog_0.wdtcnt_6_ ;
  wire watchdog_0.wdtcnt_7_ ;
  wire watchdog_0.wdtcnt_8_ ;
  wire watchdog_0.wdtcnt_9_ ;
  wire watchdog_0.wdtctl_0_ ;
  wire watchdog_0.wdtctl_1_ ;
  wire watchdog_0.wdtctl_2_ ;
  wire watchdog_0.wdtctl_3_ ;
  wire watchdog_0.wdtctl_4_ ;
  wire watchdog_0.wdtctl_5_ ;
  wire watchdog_0.wdtctl_7_ ;
  input wkup;
  INVX1 _06060_ (
    .A(multiplier_0.per_dout_0_ ),
    .Y(_00045_)
  );
  INVX1 _06061_ (
    .A(multiplier_0.per_dout_1_ ),
    .Y(_00046_)
  );
  INVX1 _06062_ (
    .A(multiplier_0.per_dout_2_ ),
    .Y(_00047_)
  );
  INVX1 _06063_ (
    .A(multiplier_0.per_dout_3_ ),
    .Y(_00000_)
  );
  INVX1 _06064_ (
    .A(multiplier_0.per_dout_4_ ),
    .Y(_00001_)
  );
  INVX1 _06065_ (
    .A(multiplier_0.per_dout_5_ ),
    .Y(_00002_)
  );
  INVX1 _06066_ (
    .A(multiplier_0.per_dout_6_ ),
    .Y(_00003_)
  );
  INVX1 _06067_ (
    .A(multiplier_0.per_dout_7_ ),
    .Y(_00004_)
  );
  INVX1 _06068_ (
    .A(multiplier_0.per_dout_8_ ),
    .Y(_00005_)
  );
  INVX1 _06069_ (
    .A(multiplier_0.per_dout_9_ ),
    .Y(_00006_)
  );
  INVX1 _06070_ (
    .A(multiplier_0.per_dout_10_ ),
    .Y(_00007_)
  );
  INVX1 _06071_ (
    .A(multiplier_0.per_dout_11_ ),
    .Y(_00008_)
  );
  INVX1 _06072_ (
    .A(multiplier_0.per_dout_12_ ),
    .Y(_00009_)
  );
  INVX1 _06073_ (
    .A(multiplier_0.per_dout_13_ ),
    .Y(_00010_)
  );
  INVX1 _06074_ (
    .A(multiplier_0.per_dout_14_ ),
    .Y(_00011_)
  );
  INVX1 _06075_ (
    .A(multiplier_0.per_dout_15_ ),
    .Y(_00012_)
  );
  NOR2X1 _06076_ (
    .A(clock_module_0.bcsctl2_rd_0_ ),
    .B(per_dout_0_),
    .Y(_00013_)
  );
  NOR2X1 _06077_ (
    .A(per_dout_sfr_0_),
    .B(per_dout_wdog_0_),
    .Y(_00014_)
  );
  NAND3X1 _06078_ (
    .A(_00045_),
    .B(_00013_),
    .C(_00014_),
    .Y(mem_backbone_0.per_dout_0_ )
  );
  NOR2X1 _06079_ (
    .A(clock_module_0.bcsctl2_rd_1_ ),
    .B(per_dout_1_),
    .Y(_00015_)
  );
  NOR2X1 _06080_ (
    .A(per_dout_sfr_1_),
    .B(per_dout_wdog_1_),
    .Y(_00016_)
  );
  NAND3X1 _06081_ (
    .A(_00046_),
    .B(_00015_),
    .C(_00016_),
    .Y(mem_backbone_0.per_dout_1_ )
  );
  NOR2X1 _06082_ (
    .A(clock_module_0.bcsctl2_rd_2_ ),
    .B(per_dout_2_),
    .Y(_00017_)
  );
  NOR2X1 _06083_ (
    .A(per_dout_sfr_2_),
    .B(per_dout_wdog_2_),
    .Y(_00018_)
  );
  NAND3X1 _06084_ (
    .A(_00047_),
    .B(_00017_),
    .C(_00018_),
    .Y(mem_backbone_0.per_dout_2_ )
  );
  NOR2X1 _06085_ (
    .A(clock_module_0.bcsctl2_rd_3_ ),
    .B(per_dout_3_),
    .Y(_00019_)
  );
  NOR2X1 _06086_ (
    .A(per_dout_sfr_3_),
    .B(per_dout_wdog_3_),
    .Y(_00020_)
  );
  NAND3X1 _06087_ (
    .A(_00000_),
    .B(_00019_),
    .C(_00020_),
    .Y(mem_backbone_0.per_dout_3_ )
  );
  NOR2X1 _06088_ (
    .A(clock_module_0.bcsctl2_rd_4_ ),
    .B(per_dout_4_),
    .Y(_00021_)
  );
  NOR2X1 _06089_ (
    .A(per_dout_sfr_4_),
    .B(per_dout_wdog_4_),
    .Y(_00022_)
  );
  NAND3X1 _06090_ (
    .A(_00001_),
    .B(_00021_),
    .C(_00022_),
    .Y(mem_backbone_0.per_dout_4_ )
  );
  NOR2X1 _06091_ (
    .A(clock_module_0.bcsctl2_rd_5_ ),
    .B(per_dout_5_),
    .Y(_00023_)
  );
  NOR2X1 _06092_ (
    .A(per_dout_sfr_5_),
    .B(per_dout_wdog_5_),
    .Y(_00024_)
  );
  NAND3X1 _06093_ (
    .A(_00002_),
    .B(_00023_),
    .C(_00024_),
    .Y(mem_backbone_0.per_dout_5_ )
  );
  NOR2X1 _06094_ (
    .A(clock_module_0.bcsctl2_rd_6_ ),
    .B(per_dout_6_),
    .Y(_00025_)
  );
  NOR2X1 _06095_ (
    .A(per_dout_sfr_6_),
    .B(per_dout_wdog_6_),
    .Y(_00026_)
  );
  NAND3X1 _06096_ (
    .A(_00003_),
    .B(_00025_),
    .C(_00026_),
    .Y(mem_backbone_0.per_dout_6_ )
  );
  NOR2X1 _06097_ (
    .A(clock_module_0.bcsctl2_rd_7_ ),
    .B(per_dout_7_),
    .Y(_00027_)
  );
  NOR2X1 _06098_ (
    .A(per_dout_sfr_7_),
    .B(per_dout_wdog_7_),
    .Y(_00028_)
  );
  NAND3X1 _06099_ (
    .A(_00004_),
    .B(_00027_),
    .C(_00028_),
    .Y(mem_backbone_0.per_dout_7_ )
  );
  NOR2X1 _06100_ (
    .A(clock_module_0.bcsctl1_rd_8_ ),
    .B(per_dout_8_),
    .Y(_00029_)
  );
  NOR2X1 _06101_ (
    .A(per_dout_sfr_8_),
    .B(per_dout_wdog_11_),
    .Y(_00030_)
  );
  NAND3X1 _06102_ (
    .A(_00005_),
    .B(_00029_),
    .C(_00030_),
    .Y(mem_backbone_0.per_dout_8_ )
  );
  NOR2X1 _06103_ (
    .A(clock_module_0.bcsctl1_rd_9_ ),
    .B(per_dout_9_),
    .Y(_00031_)
  );
  NOR2X1 _06104_ (
    .A(per_dout_sfr_9_),
    .B(1'h0),
    .Y(_00032_)
  );
  NAND3X1 _06105_ (
    .A(_00006_),
    .B(_00031_),
    .C(_00032_),
    .Y(mem_backbone_0.per_dout_9_ )
  );
  NOR2X1 _06106_ (
    .A(clock_module_0.bcsctl1_rd_10_ ),
    .B(per_dout_10_),
    .Y(_00033_)
  );
  NOR2X1 _06107_ (
    .A(per_dout_sfr_10_),
    .B(1'h0),
    .Y(_00034_)
  );
  NAND3X1 _06108_ (
    .A(_00007_),
    .B(_00033_),
    .C(_00034_),
    .Y(mem_backbone_0.per_dout_10_ )
  );
  NOR2X1 _06109_ (
    .A(clock_module_0.bcsctl1_rd_11_ ),
    .B(per_dout_11_),
    .Y(_00035_)
  );
  NOR2X1 _06110_ (
    .A(per_dout_sfr_11_),
    .B(per_dout_wdog_11_),
    .Y(_00036_)
  );
  NAND3X1 _06111_ (
    .A(_00008_),
    .B(_00035_),
    .C(_00036_),
    .Y(mem_backbone_0.per_dout_11_ )
  );
  NOR2X1 _06112_ (
    .A(clock_module_0.bcsctl1_rd_12_ ),
    .B(per_dout_12_),
    .Y(_00037_)
  );
  NOR2X1 _06113_ (
    .A(per_dout_sfr_12_),
    .B(1'h0),
    .Y(_00038_)
  );
  NAND3X1 _06114_ (
    .A(_00009_),
    .B(_00037_),
    .C(_00038_),
    .Y(mem_backbone_0.per_dout_12_ )
  );
  NOR2X1 _06115_ (
    .A(clock_module_0.bcsctl1_rd_13_ ),
    .B(per_dout_13_),
    .Y(_00039_)
  );
  NOR2X1 _06116_ (
    .A(per_dout_sfr_13_),
    .B(per_dout_wdog_11_),
    .Y(_00040_)
  );
  NAND3X1 _06117_ (
    .A(_00010_),
    .B(_00039_),
    .C(_00040_),
    .Y(mem_backbone_0.per_dout_13_ )
  );
  NOR2X1 _06118_ (
    .A(clock_module_0.bcsctl1_rd_14_ ),
    .B(per_dout_14_),
    .Y(_00041_)
  );
  NOR2X1 _06119_ (
    .A(per_dout_sfr_14_),
    .B(per_dout_wdog_11_),
    .Y(_00042_)
  );
  NAND3X1 _06120_ (
    .A(_00011_),
    .B(_00041_),
    .C(_00042_),
    .Y(mem_backbone_0.per_dout_14_ )
  );
  NOR2X1 _06121_ (
    .A(clock_module_0.bcsctl1_rd_15_ ),
    .B(per_dout_15_),
    .Y(_00043_)
  );
  NOR2X1 _06122_ (
    .A(per_dout_sfr_15_),
    .B(1'h0),
    .Y(_00044_)
  );
  NAND3X1 _06123_ (
    .A(_00012_),
    .B(_00043_),
    .C(_00044_),
    .Y(mem_backbone_0.per_dout_15_ )
  );
  BUFX2 _06124_ (
    .A(dco_clk),
    .Y(aclk)
  );
  BUFX2 _06125_ (
    .A(_00048_),
    .Y(aclk_en)
  );
  BUFX2 _06126_ (
    .A(_00049_),
    .Y(dbg_freeze)
  );
  BUFX2 _06127_ (
    .A(_00050_),
    .Y(dbg_i2c_sda_out)
  );
  BUFX2 _06128_ (
    .A(1'h1),
    .Y(dbg_uart_txd)
  );
  BUFX2 _06129_ (
    .A(1'h1),
    .Y(dco_enable)
  );
  BUFX2 _06130_ (
    .A(1'h1),
    .Y(dco_wkup)
  );
  BUFX2 _06131_ (
    .A(1'h0),
    .Y(dma_dout_0_)
  );
  BUFX2 _06132_ (
    .A(1'h0),
    .Y(dma_dout_10_)
  );
  BUFX2 _06133_ (
    .A(1'h0),
    .Y(dma_dout_11_)
  );
  BUFX2 _06134_ (
    .A(1'h0),
    .Y(dma_dout_12_)
  );
  BUFX2 _06135_ (
    .A(1'h0),
    .Y(dma_dout_13_)
  );
  BUFX2 _06136_ (
    .A(1'h0),
    .Y(dma_dout_14_)
  );
  BUFX2 _06137_ (
    .A(1'h0),
    .Y(dma_dout_15_)
  );
  BUFX2 _06138_ (
    .A(1'h0),
    .Y(dma_dout_1_)
  );
  BUFX2 _06139_ (
    .A(1'h0),
    .Y(dma_dout_2_)
  );
  BUFX2 _06140_ (
    .A(1'h0),
    .Y(dma_dout_3_)
  );
  BUFX2 _06141_ (
    .A(1'h0),
    .Y(dma_dout_4_)
  );
  BUFX2 _06142_ (
    .A(1'h0),
    .Y(dma_dout_5_)
  );
  BUFX2 _06143_ (
    .A(1'h0),
    .Y(dma_dout_6_)
  );
  BUFX2 _06144_ (
    .A(1'h0),
    .Y(dma_dout_7_)
  );
  BUFX2 _06145_ (
    .A(1'h0),
    .Y(dma_dout_8_)
  );
  BUFX2 _06146_ (
    .A(1'h0),
    .Y(dma_dout_9_)
  );
  BUFX2 _06147_ (
    .A(1'h1),
    .Y(dma_ready)
  );
  BUFX2 _06148_ (
    .A(1'h1),
    .Y(dma_resp)
  );
  BUFX2 _06149_ (
    .A(_00051_),
    .Y(dmem_addr_0_)
  );
  BUFX2 _06150_ (
    .A(_00052_),
    .Y(dmem_addr_10_)
  );
  BUFX2 _06151_ (
    .A(_00053_),
    .Y(dmem_addr_11_)
  );
  BUFX2 _06152_ (
    .A(_00054_),
    .Y(dmem_addr_12_)
  );
  BUFX2 _06153_ (
    .A(_00055_),
    .Y(dmem_addr_1_)
  );
  BUFX2 _06154_ (
    .A(_00056_),
    .Y(dmem_addr_2_)
  );
  BUFX2 _06155_ (
    .A(_00057_),
    .Y(dmem_addr_3_)
  );
  BUFX2 _06156_ (
    .A(_00058_),
    .Y(dmem_addr_4_)
  );
  BUFX2 _06157_ (
    .A(_00059_),
    .Y(dmem_addr_5_)
  );
  BUFX2 _06158_ (
    .A(_00060_),
    .Y(dmem_addr_6_)
  );
  BUFX2 _06159_ (
    .A(_00061_),
    .Y(dmem_addr_7_)
  );
  BUFX2 _06160_ (
    .A(_00062_),
    .Y(dmem_addr_8_)
  );
  BUFX2 _06161_ (
    .A(_00063_),
    .Y(dmem_addr_9_)
  );
  BUFX2 _06162_ (
    .A(_00064_),
    .Y(dmem_cen)
  );
  BUFX2 _06163_ (
    .A(_00065_),
    .Y(dmem_din_0_)
  );
  BUFX2 _06164_ (
    .A(_00066_),
    .Y(dmem_din_10_)
  );
  BUFX2 _06165_ (
    .A(_00067_),
    .Y(dmem_din_11_)
  );
  BUFX2 _06166_ (
    .A(_00068_),
    .Y(dmem_din_12_)
  );
  BUFX2 _06167_ (
    .A(_00069_),
    .Y(dmem_din_13_)
  );
  BUFX2 _06168_ (
    .A(_00070_),
    .Y(dmem_din_14_)
  );
  BUFX2 _06169_ (
    .A(_00071_),
    .Y(dmem_din_15_)
  );
  BUFX2 _06170_ (
    .A(_00072_),
    .Y(dmem_din_1_)
  );
  BUFX2 _06171_ (
    .A(_00073_),
    .Y(dmem_din_2_)
  );
  BUFX2 _06172_ (
    .A(_00074_),
    .Y(dmem_din_3_)
  );
  BUFX2 _06173_ (
    .A(_00075_),
    .Y(dmem_din_4_)
  );
  BUFX2 _06174_ (
    .A(_00076_),
    .Y(dmem_din_5_)
  );
  BUFX2 _06175_ (
    .A(_00077_),
    .Y(dmem_din_6_)
  );
  BUFX2 _06176_ (
    .A(_00078_),
    .Y(dmem_din_7_)
  );
  BUFX2 _06177_ (
    .A(_00079_),
    .Y(dmem_din_8_)
  );
  BUFX2 _06178_ (
    .A(_00080_),
    .Y(dmem_din_9_)
  );
  BUFX2 _06179_ (
    .A(_00081_),
    .Y(dmem_wen_0_)
  );
  BUFX2 _06180_ (
    .A(_00082_),
    .Y(dmem_wen_1_)
  );
  BUFX2 _06181_ (
    .A(_00083_),
    .Y(irq_acc_0_)
  );
  BUFX2 _06182_ (
    .A(_00084_),
    .Y(irq_acc_10_)
  );
  BUFX2 _06183_ (
    .A(_00085_),
    .Y(irq_acc_11_)
  );
  BUFX2 _06184_ (
    .A(_00086_),
    .Y(irq_acc_12_)
  );
  BUFX2 _06185_ (
    .A(_00087_),
    .Y(irq_acc_13_)
  );
  BUFX2 _06186_ (
    .A(_00088_),
    .Y(irq_acc_1_)
  );
  BUFX2 _06187_ (
    .A(_00089_),
    .Y(irq_acc_2_)
  );
  BUFX2 _06188_ (
    .A(_00090_),
    .Y(irq_acc_3_)
  );
  BUFX2 _06189_ (
    .A(_00091_),
    .Y(irq_acc_4_)
  );
  BUFX2 _06190_ (
    .A(_00092_),
    .Y(irq_acc_5_)
  );
  BUFX2 _06191_ (
    .A(_00093_),
    .Y(irq_acc_6_)
  );
  BUFX2 _06192_ (
    .A(_00094_),
    .Y(irq_acc_7_)
  );
  BUFX2 _06193_ (
    .A(_00095_),
    .Y(irq_acc_8_)
  );
  BUFX2 _06194_ (
    .A(_00096_),
    .Y(irq_acc_9_)
  );
  BUFX2 _06195_ (
    .A(1'h1),
    .Y(lfxt_enable)
  );
  BUFX2 _06196_ (
    .A(1'h0),
    .Y(lfxt_wkup)
  );
  BUFX2 _06197_ (
    .A(dco_clk),
    .Y(mclk)
  );
  BUFX2 _06198_ (
    .A(_00097_),
    .Y(per_addr_0_)
  );
  BUFX2 _06199_ (
    .A(_00098_),
    .Y(per_addr_10_)
  );
  BUFX2 _06200_ (
    .A(_00099_),
    .Y(per_addr_11_)
  );
  BUFX2 _06201_ (
    .A(_00100_),
    .Y(per_addr_12_)
  );
  BUFX2 _06202_ (
    .A(1'h0),
    .Y(per_addr_13_)
  );
  BUFX2 _06203_ (
    .A(_00101_),
    .Y(per_addr_1_)
  );
  BUFX2 _06204_ (
    .A(_00102_),
    .Y(per_addr_2_)
  );
  BUFX2 _06205_ (
    .A(_00103_),
    .Y(per_addr_3_)
  );
  BUFX2 _06206_ (
    .A(_00104_),
    .Y(per_addr_4_)
  );
  BUFX2 _06207_ (
    .A(_00105_),
    .Y(per_addr_5_)
  );
  BUFX2 _06208_ (
    .A(_00106_),
    .Y(per_addr_6_)
  );
  BUFX2 _06209_ (
    .A(_00107_),
    .Y(per_addr_7_)
  );
  BUFX2 _06210_ (
    .A(_00108_),
    .Y(per_addr_8_)
  );
  BUFX2 _06211_ (
    .A(_00109_),
    .Y(per_addr_9_)
  );
  BUFX2 _06212_ (
    .A(_00110_),
    .Y(per_din_0_)
  );
  BUFX2 _06213_ (
    .A(_00111_),
    .Y(per_din_10_)
  );
  BUFX2 _06214_ (
    .A(_00112_),
    .Y(per_din_11_)
  );
  BUFX2 _06215_ (
    .A(_00113_),
    .Y(per_din_12_)
  );
  BUFX2 _06216_ (
    .A(_00114_),
    .Y(per_din_13_)
  );
  BUFX2 _06217_ (
    .A(_00115_),
    .Y(per_din_14_)
  );
  BUFX2 _06218_ (
    .A(_00116_),
    .Y(per_din_15_)
  );
  BUFX2 _06219_ (
    .A(_00117_),
    .Y(per_din_1_)
  );
  BUFX2 _06220_ (
    .A(_00118_),
    .Y(per_din_2_)
  );
  BUFX2 _06221_ (
    .A(_00119_),
    .Y(per_din_3_)
  );
  BUFX2 _06222_ (
    .A(_00120_),
    .Y(per_din_4_)
  );
  BUFX2 _06223_ (
    .A(_00121_),
    .Y(per_din_5_)
  );
  BUFX2 _06224_ (
    .A(_00122_),
    .Y(per_din_6_)
  );
  BUFX2 _06225_ (
    .A(_00123_),
    .Y(per_din_7_)
  );
  BUFX2 _06226_ (
    .A(_00124_),
    .Y(per_din_8_)
  );
  BUFX2 _06227_ (
    .A(_00125_),
    .Y(per_din_9_)
  );
  BUFX2 _06228_ (
    .A(_00126_),
    .Y(per_en)
  );
  BUFX2 _06229_ (
    .A(_00127_),
    .Y(per_we_0_)
  );
  BUFX2 _06230_ (
    .A(_00128_),
    .Y(per_we_1_)
  );
  BUFX2 _06231_ (
    .A(_00129_),
    .Y(pmem_addr_0_)
  );
  BUFX2 _06232_ (
    .A(_00130_),
    .Y(pmem_addr_10_)
  );
  BUFX2 _06233_ (
    .A(_00131_),
    .Y(pmem_addr_11_)
  );
  BUFX2 _06234_ (
    .A(_00132_),
    .Y(pmem_addr_12_)
  );
  BUFX2 _06235_ (
    .A(_00133_),
    .Y(pmem_addr_13_)
  );
  BUFX2 _06236_ (
    .A(_00134_),
    .Y(pmem_addr_1_)
  );
  BUFX2 _06237_ (
    .A(_00135_),
    .Y(pmem_addr_2_)
  );
  BUFX2 _06238_ (
    .A(_00136_),
    .Y(pmem_addr_3_)
  );
  BUFX2 _06239_ (
    .A(_00137_),
    .Y(pmem_addr_4_)
  );
  BUFX2 _06240_ (
    .A(_00138_),
    .Y(pmem_addr_5_)
  );
  BUFX2 _06241_ (
    .A(_00139_),
    .Y(pmem_addr_6_)
  );
  BUFX2 _06242_ (
    .A(_00140_),
    .Y(pmem_addr_7_)
  );
  BUFX2 _06243_ (
    .A(_00141_),
    .Y(pmem_addr_8_)
  );
  BUFX2 _06244_ (
    .A(_00142_),
    .Y(pmem_addr_9_)
  );
  BUFX2 _06245_ (
    .A(_00143_),
    .Y(pmem_cen)
  );
  BUFX2 _06246_ (
    .A(_00144_),
    .Y(pmem_din_0_)
  );
  BUFX2 _06247_ (
    .A(_00145_),
    .Y(pmem_din_10_)
  );
  BUFX2 _06248_ (
    .A(_00146_),
    .Y(pmem_din_11_)
  );
  BUFX2 _06249_ (
    .A(_00147_),
    .Y(pmem_din_12_)
  );
  BUFX2 _06250_ (
    .A(_00148_),
    .Y(pmem_din_13_)
  );
  BUFX2 _06251_ (
    .A(_00149_),
    .Y(pmem_din_14_)
  );
  BUFX2 _06252_ (
    .A(_00150_),
    .Y(pmem_din_15_)
  );
  BUFX2 _06253_ (
    .A(_00151_),
    .Y(pmem_din_1_)
  );
  BUFX2 _06254_ (
    .A(_00152_),
    .Y(pmem_din_2_)
  );
  BUFX2 _06255_ (
    .A(_00153_),
    .Y(pmem_din_3_)
  );
  BUFX2 _06256_ (
    .A(_00154_),
    .Y(pmem_din_4_)
  );
  BUFX2 _06257_ (
    .A(_00155_),
    .Y(pmem_din_5_)
  );
  BUFX2 _06258_ (
    .A(_00156_),
    .Y(pmem_din_6_)
  );
  BUFX2 _06259_ (
    .A(_00157_),
    .Y(pmem_din_7_)
  );
  BUFX2 _06260_ (
    .A(_00158_),
    .Y(pmem_din_8_)
  );
  BUFX2 _06261_ (
    .A(_00159_),
    .Y(pmem_din_9_)
  );
  BUFX2 _06262_ (
    .A(_00160_),
    .Y(pmem_wen_0_)
  );
  BUFX2 _06263_ (
    .A(_00161_),
    .Y(pmem_wen_1_)
  );
  BUFX2 _06264_ (
    .A(_00162_),
    .Y(puc_rst)
  );
  BUFX2 _06265_ (
    .A(dco_clk),
    .Y(smclk)
  );
  BUFX2 _06266_ (
    .A(_00163_),
    .Y(smclk_en)
  );
  INVX1 _06267_ (
    .A(reset_n),
    .Y(clock_module_0.por_a )
  );
  INVX1 _06268_ (
    .A(_00104_),
    .Y(_00189_)
  );
  INVX1 _06269_ (
    .A(_00106_),
    .Y(_00190_)
  );
  INVX1 _06270_ (
    .A(_00100_),
    .Y(_00191_)
  );
  INVX1 _06271_ (
    .A(clock_module_0.bcsctl1_4_ ),
    .Y(_00192_)
  );
  INVX1 _06272_ (
    .A(clock_module_0.lfxt_clk_s ),
    .Y(_00193_)
  );
  INVX1 _06273_ (
    .A(clock_module_0.bcsctl2_1_ ),
    .Y(_00194_)
  );
  INVX1 _06274_ (
    .A(clock_module_0.bcsctl2_3_ ),
    .Y(_00195_)
  );
  INVX1 _06275_ (
    .A(clock_module_0.scg1 ),
    .Y(_00196_)
  );
  INVX1 _06276_ (
    .A(dbg_en),
    .Y(clock_module_0.dbg_rst_nxt )
  );
  INVX1 _06277_ (
    .A(clock_module_0.puc_noscan_n ),
    .Y(_00162_)
  );
  INVX1 _06278_ (
    .A(clock_module_0.por ),
    .Y(_00188_)
  );
  NOR2X1 _06279_ (
    .A(_00099_),
    .B(1'h0),
    .Y(_00197_)
  );
  NAND3X1 _06280_ (
    .A(_00191_),
    .B(_00126_),
    .C(_00197_),
    .Y(_00198_)
  );
  INVX1 _06281_ (
    .A(_00198_),
    .Y(_00199_)
  );
  NOR2X1 _06282_ (
    .A(_00108_),
    .B(_00107_),
    .Y(_00200_)
  );
  NOR2X1 _06283_ (
    .A(_00098_),
    .B(_00109_),
    .Y(_00201_)
  );
  NAND2X1 _06284_ (
    .A(_00200_),
    .B(_00201_),
    .Y(_00202_)
  );
  NAND2X1 _06285_ (
    .A(_00189_),
    .B(_00103_),
    .Y(_00203_)
  );
  NAND2X1 _06286_ (
    .A(_00190_),
    .B(_00105_),
    .Y(_00204_)
  );
  NOR3X1 _06287_ (
    .A(_00202_),
    .B(_00203_),
    .C(_00204_),
    .Y(_00205_)
  );
  NAND2X1 _06288_ (
    .A(_00101_),
    .B(_00097_),
    .Y(_00206_)
  );
  NOR2X1 _06289_ (
    .A(_00102_),
    .B(_00206_),
    .Y(_00207_)
  );
  NOR2X1 _06290_ (
    .A(_00108_),
    .B(_00109_),
    .Y(_00208_)
  );
  NAND3X1 _06291_ (
    .A(_00189_),
    .B(_00190_),
    .C(_00208_),
    .Y(_00209_)
  );
  NOR2X1 _06292_ (
    .A(_00107_),
    .B(_00098_),
    .Y(_00210_)
  );
  NAND3X1 _06293_ (
    .A(_00103_),
    .B(_00105_),
    .C(_00210_),
    .Y(_00211_)
  );
  NOR3X1 _06294_ (
    .A(_00198_),
    .B(_00209_),
    .C(_00211_),
    .Y(_00212_)
  );
  NAND3X1 _06295_ (
    .A(_00128_),
    .B(_00207_),
    .C(_00212_),
    .Y(_00213_)
  );
  AND2X1 _06296_ (
    .A(clock_module_0.bcsctl1_0_ ),
    .B(_00213_),
    .Y(_00168_)
  );
  AND2X1 _06297_ (
    .A(clock_module_0.bcsctl1_1_ ),
    .B(_00213_),
    .Y(_00169_)
  );
  AND2X1 _06298_ (
    .A(clock_module_0.bcsctl1_2_ ),
    .B(_00213_),
    .Y(_00170_)
  );
  AND2X1 _06299_ (
    .A(clock_module_0.bcsctl1_3_ ),
    .B(_00213_),
    .Y(_00171_)
  );
  MUX2X1 _06300_ (
    .A(clock_module_0.bcsctl1_4_ ),
    .B(_00113_),
    .S(_00213_),
    .Y(_00214_)
  );
  INVX1 _06301_ (
    .A(_00214_),
    .Y(_00172_)
  );
  MUX2X1 _06302_ (
    .A(clock_module_0.bcsctl1_5_ ),
    .B(_00114_),
    .S(_00213_),
    .Y(_00215_)
  );
  INVX1 _06303_ (
    .A(_00215_),
    .Y(_00173_)
  );
  AND2X1 _06304_ (
    .A(clock_module_0.bcsctl1_6_ ),
    .B(_00213_),
    .Y(_00174_)
  );
  AND2X1 _06305_ (
    .A(clock_module_0.bcsctl1_7_ ),
    .B(_00213_),
    .Y(_00175_)
  );
  NOR2X1 _06306_ (
    .A(clock_module_0.bcsctl1_4_ ),
    .B(clock_module_0.bcsctl1_5_ ),
    .Y(_00216_)
  );
  NAND2X1 _06307_ (
    .A(clock_module_0.bcsctl1_1_ ),
    .B(1'h1),
    .Y(_00217_)
  );
  NAND2X1 _06308_ (
    .A(clock_module_0.oscoff ),
    .B(_00217_),
    .Y(_00218_)
  );
  NOR2X1 _06309_ (
    .A(clock_module_0.lfxt_clk_dly ),
    .B(_00193_),
    .Y(_00219_)
  );
  NAND2X1 _06310_ (
    .A(_00218_),
    .B(_00219_),
    .Y(_00220_)
  );
  NOR2X1 _06311_ (
    .A(_00216_),
    .B(_00220_),
    .Y(_00221_)
  );
  NAND2X1 _06312_ (
    .A(clock_module_0.aclk_div_0_ ),
    .B(_00221_),
    .Y(_00222_)
  );
  XOR2X1 _06313_ (
    .A(clock_module_0.aclk_div_0_ ),
    .B(_00221_),
    .Y(_00164_)
  );
  NAND3X1 _06314_ (
    .A(clock_module_0.aclk_div_0_ ),
    .B(clock_module_0.aclk_div_1_ ),
    .C(_00221_),
    .Y(_00223_)
  );
  XNOR2X1 _06315_ (
    .A(clock_module_0.aclk_div_1_ ),
    .B(_00222_),
    .Y(_00165_)
  );
  XNOR2X1 _06316_ (
    .A(clock_module_0.aclk_div_2_ ),
    .B(_00223_),
    .Y(_00166_)
  );
  AOI21X1 _06317_ (
    .A(clock_module_0.bcsctl1_3_ ),
    .B(1'h1),
    .C(_00196_),
    .Y(_00224_)
  );
  AOI21X1 _06318_ (
    .A(_00218_),
    .B(_00219_),
    .C(_00195_),
    .Y(_00225_)
  );
  NOR2X1 _06319_ (
    .A(_00224_),
    .B(_00225_),
    .Y(_00226_)
  );
  NOR2X1 _06320_ (
    .A(clock_module_0.bcsctl2_1_ ),
    .B(clock_module_0.bcsctl2_2_ ),
    .Y(_00227_)
  );
  NOR3X1 _06321_ (
    .A(_00224_),
    .B(_00225_),
    .C(_00227_),
    .Y(_00228_)
  );
  AND2X1 _06322_ (
    .A(clock_module_0.smclk_div_0_ ),
    .B(_00228_),
    .Y(_00229_)
  );
  NOR2X1 _06323_ (
    .A(clock_module_0.smclk_div_0_ ),
    .B(_00228_),
    .Y(_00230_)
  );
  NOR2X1 _06324_ (
    .A(_00229_),
    .B(_00230_),
    .Y(_00184_)
  );
  NAND3X1 _06325_ (
    .A(clock_module_0.smclk_div_0_ ),
    .B(clock_module_0.smclk_div_1_ ),
    .C(_00228_),
    .Y(_00231_)
  );
  XOR2X1 _06326_ (
    .A(clock_module_0.smclk_div_1_ ),
    .B(_00229_),
    .Y(_00185_)
  );
  XNOR2X1 _06327_ (
    .A(clock_module_0.smclk_div_2_ ),
    .B(_00231_),
    .Y(_00186_)
  );
  NOR2X1 _06328_ (
    .A(_00101_),
    .B(_00097_),
    .Y(_00232_)
  );
  AND2X1 _06329_ (
    .A(_00102_),
    .B(_00232_),
    .Y(_00233_)
  );
  NAND2X1 _06330_ (
    .A(_00102_),
    .B(_00232_),
    .Y(_00234_)
  );
  NAND3X1 _06331_ (
    .A(_00127_),
    .B(_00212_),
    .C(_00233_),
    .Y(_00235_)
  );
  AND2X1 _06332_ (
    .A(clock_module_0.bcsctl2_0_ ),
    .B(_00235_),
    .Y(_00176_)
  );
  MUX2X1 _06333_ (
    .A(clock_module_0.bcsctl2_1_ ),
    .B(_00117_),
    .S(_00235_),
    .Y(_00236_)
  );
  INVX1 _06334_ (
    .A(_00236_),
    .Y(_00177_)
  );
  MUX2X1 _06335_ (
    .A(clock_module_0.bcsctl2_2_ ),
    .B(_00118_),
    .S(_00235_),
    .Y(_00237_)
  );
  INVX1 _06336_ (
    .A(_00237_),
    .Y(_00178_)
  );
  MUX2X1 _06337_ (
    .A(clock_module_0.bcsctl2_3_ ),
    .B(_00119_),
    .S(_00235_),
    .Y(_00238_)
  );
  INVX1 _06338_ (
    .A(_00238_),
    .Y(_00179_)
  );
  AND2X1 _06339_ (
    .A(clock_module_0.bcsctl2_4_ ),
    .B(_00235_),
    .Y(_00180_)
  );
  AND2X1 _06340_ (
    .A(clock_module_0.bcsctl2_5_ ),
    .B(_00235_),
    .Y(_00181_)
  );
  AND2X1 _06341_ (
    .A(clock_module_0.bcsctl2_6_ ),
    .B(_00235_),
    .Y(_00182_)
  );
  AND2X1 _06342_ (
    .A(clock_module_0.bcsctl2_7_ ),
    .B(_00235_),
    .Y(_00183_)
  );
  NOR2X1 _06343_ (
    .A(clock_module_0.dbg_rst_nxt ),
    .B(clock_module_0.puc_noscan_n ),
    .Y(_00239_)
  );
  AOI21X1 _06344_ (
    .A(clock_module_0.dbg_rst ),
    .B(_00239_),
    .C(clock_module_0.dbg_cpu_reset ),
    .Y(clock_module_0.sync_cell_puc.data_in )
  );
  NOR2X1 _06345_ (
    .A(_00128_),
    .B(_00127_),
    .Y(_00240_)
  );
  NAND3X1 _06346_ (
    .A(_00199_),
    .B(_00205_),
    .C(_00240_),
    .Y(_00241_)
  );
  NOR3X1 _06347_ (
    .A(_00102_),
    .B(_00206_),
    .C(_00241_),
    .Y(_00242_)
  );
  AND2X1 _06348_ (
    .A(clock_module_0.bcsctl1_0_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_8_ )
  );
  AND2X1 _06349_ (
    .A(clock_module_0.bcsctl1_1_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_9_ )
  );
  AND2X1 _06350_ (
    .A(clock_module_0.bcsctl1_2_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_10_ )
  );
  AND2X1 _06351_ (
    .A(clock_module_0.bcsctl1_3_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_11_ )
  );
  AND2X1 _06352_ (
    .A(clock_module_0.bcsctl1_4_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_12_ )
  );
  AND2X1 _06353_ (
    .A(clock_module_0.bcsctl1_5_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_13_ )
  );
  AND2X1 _06354_ (
    .A(clock_module_0.bcsctl1_6_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_14_ )
  );
  AND2X1 _06355_ (
    .A(clock_module_0.bcsctl1_7_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_15_ )
  );
  NOR2X1 _06356_ (
    .A(_00234_),
    .B(_00241_),
    .Y(_00243_)
  );
  AND2X1 _06357_ (
    .A(clock_module_0.bcsctl2_0_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_0_ )
  );
  AND2X1 _06358_ (
    .A(clock_module_0.bcsctl2_1_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_1_ )
  );
  AND2X1 _06359_ (
    .A(clock_module_0.bcsctl2_2_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_2_ )
  );
  AND2X1 _06360_ (
    .A(clock_module_0.bcsctl2_3_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_3_ )
  );
  AND2X1 _06361_ (
    .A(clock_module_0.bcsctl2_4_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_4_ )
  );
  AND2X1 _06362_ (
    .A(clock_module_0.bcsctl2_5_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_5_ )
  );
  AND2X1 _06363_ (
    .A(clock_module_0.bcsctl2_6_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_6_ )
  );
  AND2X1 _06364_ (
    .A(clock_module_0.bcsctl2_7_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_7_ )
  );
  OAI21X1 _06365_ (
    .A(_00192_),
    .B(clock_module_0.aclk_div_2_ ),
    .C(clock_module_0.aclk_div_1_ ),
    .Y(_00244_)
  );
  OAI21X1 _06366_ (
    .A(clock_module_0.aclk_div_0_ ),
    .B(_00216_),
    .C(cpu_en),
    .Y(_00245_)
  );
  OR2X1 _06367_ (
    .A(_00220_),
    .B(_00245_),
    .Y(_00246_)
  );
  AOI21X1 _06368_ (
    .A(clock_module_0.bcsctl1_5_ ),
    .B(_00244_),
    .C(_00246_),
    .Y(_00167_)
  );
  OAI21X1 _06369_ (
    .A(_00194_),
    .B(clock_module_0.smclk_div_2_ ),
    .C(clock_module_0.smclk_div_1_ ),
    .Y(_00247_)
  );
  OAI21X1 _06370_ (
    .A(clock_module_0.smclk_div_0_ ),
    .B(_00227_),
    .C(cpu_en),
    .Y(_00248_)
  );
  AOI21X1 _06371_ (
    .A(clock_module_0.bcsctl2_2_ ),
    .B(_00247_),
    .C(_00248_),
    .Y(_00249_)
  );
  AND2X1 _06372_ (
    .A(_00226_),
    .B(_00249_),
    .Y(_00187_)
  );
  OR2X1 _06373_ (
    .A(clock_module_0.wdt_reset ),
    .B(clock_module_0.por ),
    .Y(clock_module_0.puc_a )
  );
  DFFSR _06374_ (
    .CLK(dco_clk),
    .D(clock_module_0.dbg_rst_nxt ),
    .Q(clock_module_0.dbg_rst ),
    .R(1'h1),
    .S(_00188_)
  );
  DFFSR _06375_ (
    .CLK(dco_clk),
    .D(_00184_),
    .Q(clock_module_0.smclk_div_0_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06376_ (
    .CLK(dco_clk),
    .D(_00185_),
    .Q(clock_module_0.smclk_div_1_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06377_ (
    .CLK(dco_clk),
    .D(_00186_),
    .Q(clock_module_0.smclk_div_2_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06378_ (
    .CLK(dco_clk),
    .D(_00187_),
    .Q(_00163_),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06379_ (
    .CLK(dco_clk),
    .D(_00167_),
    .Q(_00048_),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06380_ (
    .CLK(dco_clk),
    .D(_00164_),
    .Q(clock_module_0.aclk_div_0_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06381_ (
    .CLK(dco_clk),
    .D(_00165_),
    .Q(clock_module_0.aclk_div_1_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06382_ (
    .CLK(dco_clk),
    .D(_00166_),
    .Q(clock_module_0.aclk_div_2_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06383_ (
    .CLK(dco_clk),
    .D(clock_module_0.lfxt_clk_s ),
    .Q(clock_module_0.lfxt_clk_dly ),
    .R(_00188_),
    .S(1'h1)
  );
  DFFSR _06384_ (
    .CLK(dco_clk),
    .D(_00176_),
    .Q(clock_module_0.bcsctl2_0_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06385_ (
    .CLK(dco_clk),
    .D(_00177_),
    .Q(clock_module_0.bcsctl2_1_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06386_ (
    .CLK(dco_clk),
    .D(_00178_),
    .Q(clock_module_0.bcsctl2_2_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06387_ (
    .CLK(dco_clk),
    .D(_00179_),
    .Q(clock_module_0.bcsctl2_3_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06388_ (
    .CLK(dco_clk),
    .D(_00180_),
    .Q(clock_module_0.bcsctl2_4_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06389_ (
    .CLK(dco_clk),
    .D(_00181_),
    .Q(clock_module_0.bcsctl2_5_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06390_ (
    .CLK(dco_clk),
    .D(_00182_),
    .Q(clock_module_0.bcsctl2_6_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06391_ (
    .CLK(dco_clk),
    .D(_00183_),
    .Q(clock_module_0.bcsctl2_7_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06392_ (
    .CLK(dco_clk),
    .D(_00168_),
    .Q(clock_module_0.bcsctl1_0_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06393_ (
    .CLK(dco_clk),
    .D(_00169_),
    .Q(clock_module_0.bcsctl1_1_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06394_ (
    .CLK(dco_clk),
    .D(_00170_),
    .Q(clock_module_0.bcsctl1_2_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06395_ (
    .CLK(dco_clk),
    .D(_00171_),
    .Q(clock_module_0.bcsctl1_3_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06396_ (
    .CLK(dco_clk),
    .D(_00172_),
    .Q(clock_module_0.bcsctl1_4_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06397_ (
    .CLK(dco_clk),
    .D(_00173_),
    .Q(clock_module_0.bcsctl1_5_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06398_ (
    .CLK(dco_clk),
    .D(_00174_),
    .Q(clock_module_0.bcsctl1_6_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06399_ (
    .CLK(dco_clk),
    .D(_00175_),
    .Q(clock_module_0.bcsctl1_7_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  INVX1 _06400_ (
    .A(clock_module_0.por ),
    .Y(_00250_)
  );
  DFFSR _06401_ (
    .CLK(dco_clk),
    .D(lfxt_clk),
    .Q(clock_module_0.sync_cell_lfxt_clk.data_sync_0_ ),
    .R(_00250_),
    .S(1'h1)
  );
  DFFSR _06402_ (
    .CLK(dco_clk),
    .D(clock_module_0.sync_cell_lfxt_clk.data_sync_0_ ),
    .Q(clock_module_0.lfxt_clk_s ),
    .R(_00250_),
    .S(1'h1)
  );
  INVX1 _06403_ (
    .A(clock_module_0.puc_a ),
    .Y(_00251_)
  );
  DFFSR _06404_ (
    .CLK(dco_clk),
    .D(clock_module_0.sync_cell_puc.data_in ),
    .Q(clock_module_0.sync_cell_puc.data_sync_0_ ),
    .R(_00251_),
    .S(1'h1)
  );
  DFFSR _06405_ (
    .CLK(dco_clk),
    .D(clock_module_0.sync_cell_puc.data_sync_0_ ),
    .Q(clock_module_0.puc_noscan_n ),
    .R(_00251_),
    .S(1'h1)
  );
  INVX1 _06406_ (
    .A(clock_module_0.por_a ),
    .Y(_00252_)
  );
  DFFSR _06407_ (
    .CLK(dco_clk),
    .D(1'h0),
    .Q(clock_module_0.sync_reset_por.data_sync_0_ ),
    .R(1'h1),
    .S(_00252_)
  );
  DFFSR _06408_ (
    .CLK(dco_clk),
    .D(clock_module_0.sync_reset_por.data_sync_0_ ),
    .Q(clock_module_0.por ),
    .R(1'h1),
    .S(_00252_)
  );
  INVX1 _06409_ (
    .A(dbg_0.mem_cnt_6_ ),
    .Y(_00321_)
  );
  INVX1 _06410_ (
    .A(dbg_0.mem_cnt_7_ ),
    .Y(_00322_)
  );
  INVX1 _06411_ (
    .A(dbg_0.mem_cnt_4_ ),
    .Y(_00323_)
  );
  INVX1 _06412_ (
    .A(dbg_0.mem_cnt_8_ ),
    .Y(_00324_)
  );
  INVX1 _06413_ (
    .A(dbg_0.mem_start ),
    .Y(_00325_)
  );
  INVX1 _06414_ (
    .A(dbg_0.mem_startb ),
    .Y(_00326_)
  );
  INVX1 _06415_ (
    .A(dbg_0.mem_state_0_ ),
    .Y(_00327_)
  );
  INVX1 _06416_ (
    .A(dbg_0.mem_ctl_1_ ),
    .Y(_00328_)
  );
  INVX1 _06417_ (
    .A(dbg_0.dbg_mem_addr_0_ ),
    .Y(_00329_)
  );
  INVX1 _06418_ (
    .A(dbg_0.mem_data_8_ ),
    .Y(_00330_)
  );
  INVX1 _06419_ (
    .A(dbg_0.mem_data_9_ ),
    .Y(_00331_)
  );
  INVX1 _06420_ (
    .A(dbg_0.mem_data_10_ ),
    .Y(_00332_)
  );
  INVX1 _06421_ (
    .A(dbg_0.mem_data_11_ ),
    .Y(_00333_)
  );
  INVX1 _06422_ (
    .A(dbg_0.mem_data_12_ ),
    .Y(_00334_)
  );
  INVX1 _06423_ (
    .A(dbg_0.mem_data_13_ ),
    .Y(_00335_)
  );
  INVX1 _06424_ (
    .A(dbg_0.mem_data_14_ ),
    .Y(_00336_)
  );
  INVX1 _06425_ (
    .A(dbg_0.mem_data_15_ ),
    .Y(_00337_)
  );
  INVX1 _06426_ (
    .A(dbg_0.dbg_rd_rdy ),
    .Y(_00338_)
  );
  INVX1 _06427_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00339_)
  );
  INVX1 _06428_ (
    .A(dbg_0.dbg_addr_0_ ),
    .Y(_00340_)
  );
  INVX1 _06429_ (
    .A(dbg_0.dbg_mem_addr_1_ ),
    .Y(_00341_)
  );
  INVX1 _06430_ (
    .A(dbg_0.dbg_mem_addr_2_ ),
    .Y(_00342_)
  );
  INVX1 _06431_ (
    .A(dbg_0.dbg_din_2_ ),
    .Y(_00343_)
  );
  INVX1 _06432_ (
    .A(dbg_0.dbg_mem_addr_3_ ),
    .Y(_00344_)
  );
  INVX1 _06433_ (
    .A(dbg_0.dbg_din_3_ ),
    .Y(_00345_)
  );
  INVX1 _06434_ (
    .A(dbg_0.dbg_mem_addr_4_ ),
    .Y(_00346_)
  );
  INVX1 _06435_ (
    .A(dbg_0.dbg_mem_addr_5_ ),
    .Y(_00347_)
  );
  INVX1 _06436_ (
    .A(dbg_0.dbg_mem_addr_6_ ),
    .Y(_00348_)
  );
  INVX1 _06437_ (
    .A(dbg_0.dbg_din_6_ ),
    .Y(_00349_)
  );
  INVX1 _06438_ (
    .A(dbg_0.dbg_mem_addr_7_ ),
    .Y(_00350_)
  );
  INVX1 _06439_ (
    .A(dbg_0.dbg_din_7_ ),
    .Y(_00351_)
  );
  INVX1 _06440_ (
    .A(dbg_0.dbg_mem_addr_8_ ),
    .Y(_00352_)
  );
  INVX1 _06441_ (
    .A(dbg_0.dbg_din_8_ ),
    .Y(_00353_)
  );
  INVX1 _06442_ (
    .A(dbg_0.dbg_mem_addr_9_ ),
    .Y(_00354_)
  );
  INVX1 _06443_ (
    .A(dbg_0.dbg_mem_addr_10_ ),
    .Y(_00355_)
  );
  INVX1 _06444_ (
    .A(dbg_0.dbg_mem_addr_11_ ),
    .Y(_00356_)
  );
  INVX1 _06445_ (
    .A(dbg_0.dbg_din_11_ ),
    .Y(_00357_)
  );
  INVX1 _06446_ (
    .A(dbg_0.dbg_mem_addr_12_ ),
    .Y(_00358_)
  );
  INVX1 _06447_ (
    .A(dbg_0.dbg_din_12_ ),
    .Y(_00359_)
  );
  INVX1 _06448_ (
    .A(dbg_0.dbg_din_14_ ),
    .Y(_00360_)
  );
  INVX1 _06449_ (
    .A(dbg_0.dbg_mem_rd_dly ),
    .Y(_00361_)
  );
  INVX1 _06450_ (
    .A(dbg_0.fe_mdb_in_6_ ),
    .Y(_00362_)
  );
  INVX1 _06451_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .Y(_00363_)
  );
  INVX1 _06452_ (
    .A(cpu_en),
    .Y(_00364_)
  );
  INVX1 _06453_ (
    .A(clock_module_0.dbg_rst ),
    .Y(_00320_)
  );
  NOR2X1 _06454_ (
    .A(dbg_0.mem_cnt_0_ ),
    .B(dbg_0.mem_cnt_1_ ),
    .Y(_00365_)
  );
  NOR2X1 _06455_ (
    .A(dbg_0.mem_cnt_2_ ),
    .B(dbg_0.mem_cnt_3_ ),
    .Y(_00366_)
  );
  AND2X1 _06456_ (
    .A(_00365_),
    .B(_00366_),
    .Y(_00367_)
  );
  NAND2X1 _06457_ (
    .A(_00365_),
    .B(_00366_),
    .Y(_00368_)
  );
  NOR2X1 _06458_ (
    .A(dbg_0.mem_cnt_14_ ),
    .B(dbg_0.mem_cnt_15_ ),
    .Y(_00369_)
  );
  OR2X1 _06459_ (
    .A(dbg_0.mem_cnt_14_ ),
    .B(dbg_0.mem_cnt_15_ ),
    .Y(_00370_)
  );
  NOR2X1 _06460_ (
    .A(dbg_0.mem_cnt_12_ ),
    .B(dbg_0.mem_cnt_13_ ),
    .Y(_00371_)
  );
  OR2X1 _06461_ (
    .A(dbg_0.mem_cnt_12_ ),
    .B(dbg_0.mem_cnt_13_ ),
    .Y(_00372_)
  );
  NOR2X1 _06462_ (
    .A(dbg_0.mem_cnt_8_ ),
    .B(dbg_0.mem_cnt_9_ ),
    .Y(_00373_)
  );
  OR2X1 _06463_ (
    .A(dbg_0.mem_cnt_8_ ),
    .B(dbg_0.mem_cnt_9_ ),
    .Y(_00374_)
  );
  NOR2X1 _06464_ (
    .A(dbg_0.mem_cnt_10_ ),
    .B(dbg_0.mem_cnt_11_ ),
    .Y(_00375_)
  );
  OR2X1 _06465_ (
    .A(dbg_0.mem_cnt_10_ ),
    .B(dbg_0.mem_cnt_11_ ),
    .Y(_00376_)
  );
  NOR2X1 _06466_ (
    .A(dbg_0.mem_cnt_4_ ),
    .B(dbg_0.mem_cnt_5_ ),
    .Y(_00377_)
  );
  OR2X1 _06467_ (
    .A(dbg_0.mem_cnt_4_ ),
    .B(dbg_0.mem_cnt_5_ ),
    .Y(_00378_)
  );
  NOR2X1 _06468_ (
    .A(dbg_0.mem_cnt_6_ ),
    .B(dbg_0.mem_cnt_7_ ),
    .Y(_00379_)
  );
  OR2X1 _06469_ (
    .A(dbg_0.mem_cnt_6_ ),
    .B(dbg_0.mem_cnt_7_ ),
    .Y(_00380_)
  );
  NOR3X1 _06470_ (
    .A(_00370_),
    .B(_00374_),
    .C(_00376_),
    .Y(_00381_)
  );
  NAND3X1 _06471_ (
    .A(_00369_),
    .B(_00373_),
    .C(_00375_),
    .Y(_00382_)
  );
  NOR3X1 _06472_ (
    .A(_00372_),
    .B(_00378_),
    .C(_00380_),
    .Y(_00383_)
  );
  NAND3X1 _06473_ (
    .A(_00371_),
    .B(_00377_),
    .C(_00379_),
    .Y(_00384_)
  );
  NOR3X1 _06474_ (
    .A(_00368_),
    .B(_00382_),
    .C(_00384_),
    .Y(_00385_)
  );
  NAND3X1 _06475_ (
    .A(_00367_),
    .B(_00381_),
    .C(_00383_),
    .Y(_00386_)
  );
  OAI21X1 _06476_ (
    .A(_00325_),
    .B(_00386_),
    .C(_00326_),
    .Y(_00387_)
  );
  NOR2X1 _06477_ (
    .A(dbg_0.mem_state_1_ ),
    .B(dbg_0.mem_state_3_ ),
    .Y(_00388_)
  );
  OAI21X1 _06478_ (
    .A(_00327_),
    .B(_00387_),
    .C(_00388_),
    .Y(_00318_)
  );
  NOR2X1 _06479_ (
    .A(dbg_0.mem_ctl_2_ ),
    .B(_00388_),
    .Y(dbg_0.dbg_mem_en )
  );
  OAI21X1 _06480_ (
    .A(dbg_0.mem_state_1_ ),
    .B(dbg_0.mem_state_3_ ),
    .C(dbg_0.mem_ctl_1_ ),
    .Y(_00389_)
  );
  INVX1 _06481_ (
    .A(_00389_),
    .Y(_00390_)
  );
  NAND2X1 _06482_ (
    .A(dbg_0.mem_ctl_1_ ),
    .B(dbg_0.dbg_mem_en ),
    .Y(_00391_)
  );
  AOI21X1 _06483_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00329_),
    .C(_00391_),
    .Y(dbg_0.dbg_mem_wr_1_ )
  );
  AND2X1 _06484_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(dbg_0.dbg_mem_addr_0_ ),
    .Y(_00392_)
  );
  NAND2X1 _06485_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(dbg_0.dbg_mem_addr_0_ ),
    .Y(_00393_)
  );
  NOR2X1 _06486_ (
    .A(_00391_),
    .B(_00392_),
    .Y(dbg_0.dbg_mem_wr_0_ )
  );
  AND2X1 _06487_ (
    .A(dbg_0.mem_state_0_ ),
    .B(_00387_),
    .Y(_00394_)
  );
  AND2X1 _06488_ (
    .A(cpu_halt_st),
    .B(_00394_),
    .Y(_00317_)
  );
  AND2X1 _06489_ (
    .A(cpu_halt_st),
    .B(dbg_0.mem_state_2_ ),
    .Y(_00316_)
  );
  NOR2X1 _06490_ (
    .A(dbg_0.mem_state_2_ ),
    .B(_00394_),
    .Y(_00395_)
  );
  NOR2X1 _06491_ (
    .A(cpu_halt_st),
    .B(_00395_),
    .Y(_00319_)
  );
  AND2X1 _06492_ (
    .A(dbg_0.mem_data_0_ ),
    .B(_00393_),
    .Y(_00144_)
  );
  AND2X1 _06493_ (
    .A(dbg_0.mem_data_1_ ),
    .B(_00393_),
    .Y(_00151_)
  );
  AND2X1 _06494_ (
    .A(dbg_0.mem_data_2_ ),
    .B(_00393_),
    .Y(_00152_)
  );
  AND2X1 _06495_ (
    .A(dbg_0.mem_data_3_ ),
    .B(_00393_),
    .Y(_00153_)
  );
  AND2X1 _06496_ (
    .A(dbg_0.mem_data_4_ ),
    .B(_00393_),
    .Y(_00154_)
  );
  AND2X1 _06497_ (
    .A(dbg_0.mem_data_5_ ),
    .B(_00393_),
    .Y(_00155_)
  );
  AND2X1 _06498_ (
    .A(dbg_0.mem_data_6_ ),
    .B(_00393_),
    .Y(_00156_)
  );
  AND2X1 _06499_ (
    .A(dbg_0.mem_data_7_ ),
    .B(_00393_),
    .Y(_00157_)
  );
  NAND2X1 _06500_ (
    .A(dbg_0.mem_data_0_ ),
    .B(_00392_),
    .Y(_00396_)
  );
  OAI21X1 _06501_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00330_),
    .C(_00396_),
    .Y(_00158_)
  );
  NAND2X1 _06502_ (
    .A(dbg_0.mem_data_1_ ),
    .B(_00392_),
    .Y(_00397_)
  );
  OAI21X1 _06503_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00331_),
    .C(_00397_),
    .Y(_00159_)
  );
  NAND2X1 _06504_ (
    .A(dbg_0.mem_data_2_ ),
    .B(_00392_),
    .Y(_00398_)
  );
  OAI21X1 _06505_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00332_),
    .C(_00398_),
    .Y(_00145_)
  );
  NAND2X1 _06506_ (
    .A(dbg_0.mem_data_3_ ),
    .B(_00392_),
    .Y(_00399_)
  );
  OAI21X1 _06507_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00333_),
    .C(_00399_),
    .Y(_00146_)
  );
  NAND2X1 _06508_ (
    .A(dbg_0.mem_data_4_ ),
    .B(_00392_),
    .Y(_00400_)
  );
  OAI21X1 _06509_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00334_),
    .C(_00400_),
    .Y(_00147_)
  );
  NAND2X1 _06510_ (
    .A(dbg_0.mem_data_5_ ),
    .B(_00392_),
    .Y(_00401_)
  );
  OAI21X1 _06511_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00335_),
    .C(_00401_),
    .Y(_00148_)
  );
  NAND2X1 _06512_ (
    .A(dbg_0.mem_data_6_ ),
    .B(_00392_),
    .Y(_00402_)
  );
  OAI21X1 _06513_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00336_),
    .C(_00402_),
    .Y(_00149_)
  );
  NAND2X1 _06514_ (
    .A(dbg_0.mem_data_7_ ),
    .B(_00392_),
    .Y(_00403_)
  );
  OAI21X1 _06515_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00337_),
    .C(_00403_),
    .Y(_00150_)
  );
  NOR2X1 _06516_ (
    .A(dbg_0.dbg_rd_rdy ),
    .B(dbg_0.dbg_i2c_0.dbg_wr ),
    .Y(_00404_)
  );
  NOR2X1 _06517_ (
    .A(_00386_),
    .B(_00404_),
    .Y(dbg_0.dbg_i2c_0.mem_burst_end )
  );
  AOI21X1 _06518_ (
    .A(_00338_),
    .B(_00389_),
    .C(_00339_),
    .Y(_00405_)
  );
  OAI21X1 _06519_ (
    .A(dbg_0.dbg_rd_rdy ),
    .B(_00390_),
    .C(dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00406_)
  );
  NOR2X1 _06520_ (
    .A(_00385_),
    .B(_00406_),
    .Y(_00407_)
  );
  NAND2X1 _06521_ (
    .A(_00386_),
    .B(_00405_),
    .Y(_00408_)
  );
  OR2X1 _06522_ (
    .A(dbg_0.mem_ctl_2_ ),
    .B(dbg_0.dbg_i2c_0.mem_bw ),
    .Y(_00409_)
  );
  NAND3X1 _06523_ (
    .A(_00386_),
    .B(_00405_),
    .C(_00409_),
    .Y(_00410_)
  );
  OR2X1 _06524_ (
    .A(_00329_),
    .B(_00410_),
    .Y(_00411_)
  );
  XNOR2X1 _06525_ (
    .A(dbg_0.dbg_mem_addr_0_ ),
    .B(_00410_),
    .Y(_00412_)
  );
  NOR2X1 _06526_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_addr_1_ ),
    .Y(_00413_)
  );
  NAND2X1 _06527_ (
    .A(dbg_0.dbg_addr_0_ ),
    .B(_00413_),
    .Y(_00414_)
  );
  OR2X1 _06528_ (
    .A(dbg_0.dbg_addr_3_ ),
    .B(dbg_0.dbg_addr_4_ ),
    .Y(_00415_)
  );
  NOR2X1 _06529_ (
    .A(dbg_0.dbg_addr_5_ ),
    .B(_00415_),
    .Y(_00416_)
  );
  NAND2X1 _06530_ (
    .A(dbg_0.dbg_addr_2_ ),
    .B(_00416_),
    .Y(_00417_)
  );
  NOR2X1 _06531_ (
    .A(_00414_),
    .B(_00417_),
    .Y(_00418_)
  );
  NAND2X1 _06532_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00418_),
    .Y(_00419_)
  );
  NOR2X1 _06533_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_addr_2_ ),
    .Y(_00420_)
  );
  AOI21X1 _06534_ (
    .A(dbg_0.dbg_addr_2_ ),
    .B(_00416_),
    .C(dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00421_)
  );
  NOR2X1 _06535_ (
    .A(_00414_),
    .B(_00421_),
    .Y(_00422_)
  );
  AND2X1 _06536_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00422_),
    .Y(_00423_)
  );
  NAND2X1 _06537_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00422_),
    .Y(_00424_)
  );
  MUX2X1 _06538_ (
    .A(dbg_0.dbg_din_0_ ),
    .B(_00412_),
    .S(_00423_),
    .Y(_00425_)
  );
  INVX1 _06539_ (
    .A(_00425_),
    .Y(_00262_)
  );
  NOR2X1 _06540_ (
    .A(_00408_),
    .B(_00409_),
    .Y(_00426_)
  );
  NOR3X1 _06541_ (
    .A(_00341_),
    .B(_00408_),
    .C(_00409_),
    .Y(_00427_)
  );
  NOR2X1 _06542_ (
    .A(dbg_0.dbg_mem_addr_1_ ),
    .B(_00426_),
    .Y(_00428_)
  );
  OAI21X1 _06543_ (
    .A(_00427_),
    .B(_00428_),
    .C(_00411_),
    .Y(_00429_)
  );
  NOR3X1 _06544_ (
    .A(_00329_),
    .B(_00341_),
    .C(_00410_),
    .Y(_00430_)
  );
  OAI21X1 _06545_ (
    .A(_00341_),
    .B(_00411_),
    .C(_00429_),
    .Y(_00431_)
  );
  NAND2X1 _06546_ (
    .A(dbg_0.dbg_din_1_ ),
    .B(_00423_),
    .Y(_00432_)
  );
  OAI21X1 _06547_ (
    .A(_00423_),
    .B(_00431_),
    .C(_00432_),
    .Y(_00269_)
  );
  NOR2X1 _06548_ (
    .A(_00427_),
    .B(_00430_),
    .Y(_00433_)
  );
  NOR2X1 _06549_ (
    .A(_00342_),
    .B(_00433_),
    .Y(_00434_)
  );
  OAI21X1 _06550_ (
    .A(_00427_),
    .B(_00430_),
    .C(dbg_0.dbg_mem_addr_2_ ),
    .Y(_00435_)
  );
  NAND2X1 _06551_ (
    .A(_00342_),
    .B(_00433_),
    .Y(_00436_)
  );
  NAND3X1 _06552_ (
    .A(_00424_),
    .B(_00435_),
    .C(_00436_),
    .Y(_00437_)
  );
  OAI21X1 _06553_ (
    .A(_00343_),
    .B(_00424_),
    .C(_00437_),
    .Y(_00270_)
  );
  NOR2X1 _06554_ (
    .A(_00344_),
    .B(_00435_),
    .Y(_00438_)
  );
  OAI21X1 _06555_ (
    .A(dbg_0.dbg_mem_addr_3_ ),
    .B(_00434_),
    .C(_00419_),
    .Y(_00439_)
  );
  OAI22X1 _06556_ (
    .A(_00345_),
    .B(_00424_),
    .C(_00438_),
    .D(_00439_),
    .Y(_00271_)
  );
  OAI21X1 _06557_ (
    .A(_00344_),
    .B(_00435_),
    .C(_00346_),
    .Y(_00440_)
  );
  NOR3X1 _06558_ (
    .A(_00344_),
    .B(_00346_),
    .C(_00435_),
    .Y(_00441_)
  );
  NAND3X1 _06559_ (
    .A(dbg_0.dbg_mem_addr_3_ ),
    .B(dbg_0.dbg_mem_addr_4_ ),
    .C(_00434_),
    .Y(_00442_)
  );
  NAND2X1 _06560_ (
    .A(_00440_),
    .B(_00442_),
    .Y(_00443_)
  );
  NAND2X1 _06561_ (
    .A(dbg_0.dbg_din_4_ ),
    .B(_00423_),
    .Y(_00444_)
  );
  OAI21X1 _06562_ (
    .A(_00423_),
    .B(_00443_),
    .C(_00444_),
    .Y(_00272_)
  );
  NOR2X1 _06563_ (
    .A(dbg_0.dbg_mem_addr_5_ ),
    .B(_00441_),
    .Y(_00445_)
  );
  OAI21X1 _06564_ (
    .A(_00347_),
    .B(_00442_),
    .C(_00419_),
    .Y(_00446_)
  );
  NAND2X1 _06565_ (
    .A(dbg_0.dbg_din_5_ ),
    .B(_00423_),
    .Y(_00447_)
  );
  OAI21X1 _06566_ (
    .A(_00445_),
    .B(_00446_),
    .C(_00447_),
    .Y(_00273_)
  );
  NAND3X1 _06567_ (
    .A(dbg_0.dbg_mem_addr_5_ ),
    .B(dbg_0.dbg_mem_addr_6_ ),
    .C(_00441_),
    .Y(_00448_)
  );
  OAI21X1 _06568_ (
    .A(_00347_),
    .B(_00442_),
    .C(_00348_),
    .Y(_00449_)
  );
  NAND2X1 _06569_ (
    .A(_00448_),
    .B(_00449_),
    .Y(_00450_)
  );
  NAND2X1 _06570_ (
    .A(dbg_0.dbg_din_6_ ),
    .B(_00423_),
    .Y(_00451_)
  );
  OAI21X1 _06571_ (
    .A(_00423_),
    .B(_00450_),
    .C(_00451_),
    .Y(_00274_)
  );
  NOR2X1 _06572_ (
    .A(_00350_),
    .B(_00448_),
    .Y(_00452_)
  );
  XNOR2X1 _06573_ (
    .A(_00350_),
    .B(_00448_),
    .Y(_00453_)
  );
  NAND2X1 _06574_ (
    .A(dbg_0.dbg_din_7_ ),
    .B(_00423_),
    .Y(_00454_)
  );
  OAI21X1 _06575_ (
    .A(_00423_),
    .B(_00453_),
    .C(_00454_),
    .Y(_00275_)
  );
  NOR3X1 _06576_ (
    .A(_00350_),
    .B(_00352_),
    .C(_00448_),
    .Y(_00455_)
  );
  NAND2X1 _06577_ (
    .A(dbg_0.dbg_mem_addr_8_ ),
    .B(_00452_),
    .Y(_00456_)
  );
  OAI21X1 _06578_ (
    .A(dbg_0.dbg_mem_addr_8_ ),
    .B(_00452_),
    .C(_00419_),
    .Y(_00457_)
  );
  OAI22X1 _06579_ (
    .A(_00353_),
    .B(_00424_),
    .C(_00455_),
    .D(_00457_),
    .Y(_00276_)
  );
  XNOR2X1 _06580_ (
    .A(dbg_0.dbg_mem_addr_9_ ),
    .B(_00455_),
    .Y(_00458_)
  );
  NAND2X1 _06581_ (
    .A(dbg_0.dbg_din_9_ ),
    .B(_00423_),
    .Y(_00459_)
  );
  OAI21X1 _06582_ (
    .A(_00423_),
    .B(_00458_),
    .C(_00459_),
    .Y(_00277_)
  );
  NAND3X1 _06583_ (
    .A(dbg_0.dbg_mem_addr_9_ ),
    .B(dbg_0.dbg_mem_addr_10_ ),
    .C(_00455_),
    .Y(_00460_)
  );
  OAI21X1 _06584_ (
    .A(_00354_),
    .B(_00456_),
    .C(_00355_),
    .Y(_00461_)
  );
  NAND2X1 _06585_ (
    .A(_00460_),
    .B(_00461_),
    .Y(_00462_)
  );
  NAND2X1 _06586_ (
    .A(dbg_0.dbg_din_10_ ),
    .B(_00423_),
    .Y(_00463_)
  );
  OAI21X1 _06587_ (
    .A(_00423_),
    .B(_00462_),
    .C(_00463_),
    .Y(_00263_)
  );
  XNOR2X1 _06588_ (
    .A(_00356_),
    .B(_00460_),
    .Y(_00464_)
  );
  NAND2X1 _06589_ (
    .A(dbg_0.dbg_din_11_ ),
    .B(_00423_),
    .Y(_00465_)
  );
  OAI21X1 _06590_ (
    .A(_00423_),
    .B(_00464_),
    .C(_00465_),
    .Y(_00264_)
  );
  NOR3X1 _06591_ (
    .A(_00356_),
    .B(_00358_),
    .C(_00460_),
    .Y(_00466_)
  );
  OAI21X1 _06592_ (
    .A(_00356_),
    .B(_00460_),
    .C(_00358_),
    .Y(_00467_)
  );
  NAND2X1 _06593_ (
    .A(_00419_),
    .B(_00467_),
    .Y(_00468_)
  );
  OAI22X1 _06594_ (
    .A(_00359_),
    .B(_00424_),
    .C(_00466_),
    .D(_00468_),
    .Y(_00265_)
  );
  NAND2X1 _06595_ (
    .A(dbg_0.dbg_mem_addr_13_ ),
    .B(_00466_),
    .Y(_00469_)
  );
  XNOR2X1 _06596_ (
    .A(dbg_0.dbg_mem_addr_13_ ),
    .B(_00466_),
    .Y(_00470_)
  );
  NAND2X1 _06597_ (
    .A(dbg_0.dbg_din_13_ ),
    .B(_00423_),
    .Y(_00471_)
  );
  OAI21X1 _06598_ (
    .A(_00423_),
    .B(_00470_),
    .C(_00471_),
    .Y(_00266_)
  );
  NAND3X1 _06599_ (
    .A(dbg_0.dbg_mem_addr_13_ ),
    .B(dbg_0.dbg_mem_addr_14_ ),
    .C(_00466_),
    .Y(_00472_)
  );
  XOR2X1 _06600_ (
    .A(dbg_0.dbg_mem_addr_14_ ),
    .B(_00469_),
    .Y(_00473_)
  );
  NAND2X1 _06601_ (
    .A(dbg_0.dbg_din_14_ ),
    .B(_00423_),
    .Y(_00474_)
  );
  OAI21X1 _06602_ (
    .A(_00423_),
    .B(_00473_),
    .C(_00474_),
    .Y(_00267_)
  );
  XOR2X1 _06603_ (
    .A(dbg_0.dbg_mem_addr_15_ ),
    .B(_00472_),
    .Y(_00475_)
  );
  NOR2X1 _06604_ (
    .A(dbg_0.dbg_din_15_ ),
    .B(_00424_),
    .Y(_00476_)
  );
  AOI21X1 _06605_ (
    .A(_00424_),
    .B(_00475_),
    .C(_00476_),
    .Y(_00268_)
  );
  NAND2X1 _06606_ (
    .A(dbg_0.mem_start ),
    .B(_00386_),
    .Y(_00477_)
  );
  NOR2X1 _06607_ (
    .A(dbg_0.mem_ctl_1_ ),
    .B(_00477_),
    .Y(dbg_0.dbg_i2c_0.mem_burst_rd )
  );
  NOR2X1 _06608_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_i2c_0.mem_burst_rd ),
    .Y(_00478_)
  );
  OAI21X1 _06609_ (
    .A(dbg_0.mem_state_1_ ),
    .B(dbg_0.mem_state_3_ ),
    .C(dbg_0.mem_ctl_2_ ),
    .Y(_00479_)
  );
  NOR2X1 _06610_ (
    .A(dbg_0.mem_ctl_1_ ),
    .B(_00479_),
    .Y(_00480_)
  );
  NOR2X1 _06611_ (
    .A(dbg_0.dbg_mem_rd_dly ),
    .B(_00480_),
    .Y(_00481_)
  );
  NAND2X1 _06612_ (
    .A(dbg_0.dbg_i2c_0.dbg_rd ),
    .B(_00478_),
    .Y(_00482_)
  );
  OAI21X1 _06613_ (
    .A(_00478_),
    .B(_00481_),
    .C(_00482_),
    .Y(_00259_)
  );
  AOI21X1 _06614_ (
    .A(_00340_),
    .B(dbg_0.dbg_addr_1_ ),
    .C(dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00483_)
  );
  NAND2X1 _06615_ (
    .A(_00416_),
    .B(_00420_),
    .Y(_00484_)
  );
  NOR2X1 _06616_ (
    .A(_00483_),
    .B(_00484_),
    .Y(_00485_)
  );
  AND2X1 _06617_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00485_),
    .Y(_00486_)
  );
  NAND3X1 _06618_ (
    .A(cpu_halt_st),
    .B(dbg_0.dbg_din_2_ ),
    .C(_00486_),
    .Y(_00487_)
  );
  INVX1 _06619_ (
    .A(_00487_),
    .Y(dbg_0.istep )
  );
  OR2X1 _06620_ (
    .A(dbg_0.inc_step_0_ ),
    .B(dbg_0.istep ),
    .Y(_00261_)
  );
  NAND3X1 _06621_ (
    .A(_00339_),
    .B(dbg_0.dbg_addr_0_ ),
    .C(dbg_0.dbg_addr_1_ ),
    .Y(_00488_)
  );
  NOR2X1 _06622_ (
    .A(_00421_),
    .B(_00488_),
    .Y(_00489_)
  );
  AND2X1 _06623_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00489_),
    .Y(_00490_)
  );
  NAND2X1 _06624_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00489_),
    .Y(_00491_)
  );
  OR2X1 _06625_ (
    .A(dbg_0.mem_cnt_0_ ),
    .B(_00408_),
    .Y(_00492_)
  );
  OAI21X1 _06626_ (
    .A(_00385_),
    .B(_00406_),
    .C(dbg_0.mem_cnt_0_ ),
    .Y(_00493_)
  );
  AND2X1 _06627_ (
    .A(_00492_),
    .B(_00493_),
    .Y(_00494_)
  );
  NAND2X1 _06628_ (
    .A(dbg_0.dbg_din_0_ ),
    .B(_00490_),
    .Y(_00495_)
  );
  OAI21X1 _06629_ (
    .A(_00490_),
    .B(_00494_),
    .C(_00495_),
    .Y(_00279_)
  );
  OR2X1 _06630_ (
    .A(dbg_0.mem_cnt_1_ ),
    .B(_00492_),
    .Y(_00496_)
  );
  OAI21X1 _06631_ (
    .A(dbg_0.mem_cnt_0_ ),
    .B(_00408_),
    .C(dbg_0.mem_cnt_1_ ),
    .Y(_00497_)
  );
  AND2X1 _06632_ (
    .A(_00496_),
    .B(_00497_),
    .Y(_00498_)
  );
  NAND2X1 _06633_ (
    .A(dbg_0.dbg_din_1_ ),
    .B(_00490_),
    .Y(_00499_)
  );
  OAI21X1 _06634_ (
    .A(_00490_),
    .B(_00498_),
    .C(_00499_),
    .Y(_00286_)
  );
  NOR2X1 _06635_ (
    .A(dbg_0.mem_cnt_2_ ),
    .B(_00496_),
    .Y(_00500_)
  );
  AND2X1 _06636_ (
    .A(dbg_0.mem_cnt_2_ ),
    .B(_00496_),
    .Y(_00501_)
  );
  OAI21X1 _06637_ (
    .A(_00500_),
    .B(_00501_),
    .C(_00491_),
    .Y(_00502_)
  );
  OAI21X1 _06638_ (
    .A(_00343_),
    .B(_00491_),
    .C(_00502_),
    .Y(_00287_)
  );
  XNOR2X1 _06639_ (
    .A(dbg_0.mem_cnt_3_ ),
    .B(_00500_),
    .Y(_00503_)
  );
  NAND2X1 _06640_ (
    .A(dbg_0.dbg_din_3_ ),
    .B(_00490_),
    .Y(_00504_)
  );
  OAI21X1 _06641_ (
    .A(_00490_),
    .B(_00503_),
    .C(_00504_),
    .Y(_00288_)
  );
  NAND2X1 _06642_ (
    .A(dbg_0.mem_cnt_4_ ),
    .B(_00407_),
    .Y(_00505_)
  );
  NAND2X1 _06643_ (
    .A(_00368_),
    .B(_00405_),
    .Y(_00506_)
  );
  NOR2X1 _06644_ (
    .A(dbg_0.mem_cnt_4_ ),
    .B(_00506_),
    .Y(_00507_)
  );
  AOI21X1 _06645_ (
    .A(_00323_),
    .B(_00408_),
    .C(_00507_),
    .Y(_00508_)
  );
  OAI21X1 _06646_ (
    .A(_00368_),
    .B(_00505_),
    .C(_00508_),
    .Y(_00509_)
  );
  NAND2X1 _06647_ (
    .A(dbg_0.dbg_din_4_ ),
    .B(_00490_),
    .Y(_00510_)
  );
  OAI21X1 _06648_ (
    .A(_00490_),
    .B(_00509_),
    .C(_00510_),
    .Y(_00289_)
  );
  NOR2X1 _06649_ (
    .A(dbg_0.dbg_din_5_ ),
    .B(_00491_),
    .Y(_00511_)
  );
  OAI21X1 _06650_ (
    .A(_00323_),
    .B(_00408_),
    .C(_00506_),
    .Y(_00512_)
  );
  XNOR2X1 _06651_ (
    .A(dbg_0.mem_cnt_5_ ),
    .B(_00407_),
    .Y(_00513_)
  );
  XOR2X1 _06652_ (
    .A(_00512_),
    .B(_00513_),
    .Y(_00514_)
  );
  AOI21X1 _06653_ (
    .A(_00491_),
    .B(_00514_),
    .C(_00511_),
    .Y(_00290_)
  );
  OAI21X1 _06654_ (
    .A(_00368_),
    .B(_00378_),
    .C(_00407_),
    .Y(_00515_)
  );
  XNOR2X1 _06655_ (
    .A(dbg_0.mem_cnt_6_ ),
    .B(_00407_),
    .Y(_00516_)
  );
  MUX2X1 _06656_ (
    .A(_00516_),
    .B(_00321_),
    .S(_00515_),
    .Y(_00517_)
  );
  NAND2X1 _06657_ (
    .A(_00491_),
    .B(_00517_),
    .Y(_00518_)
  );
  OAI21X1 _06658_ (
    .A(_00349_),
    .B(_00491_),
    .C(_00518_),
    .Y(_00291_)
  );
  OAI21X1 _06659_ (
    .A(_00321_),
    .B(_00408_),
    .C(_00515_),
    .Y(_00519_)
  );
  OAI21X1 _06660_ (
    .A(_00385_),
    .B(_00406_),
    .C(_00322_),
    .Y(_00520_)
  );
  NAND3X1 _06661_ (
    .A(dbg_0.mem_cnt_7_ ),
    .B(_00386_),
    .C(_00405_),
    .Y(_00521_)
  );
  AND2X1 _06662_ (
    .A(_00520_),
    .B(_00521_),
    .Y(_00522_)
  );
  MUX2X1 _06663_ (
    .A(dbg_0.mem_cnt_7_ ),
    .B(_00522_),
    .S(_00519_),
    .Y(_00523_)
  );
  MUX2X1 _06664_ (
    .A(_00351_),
    .B(_00523_),
    .S(_00490_),
    .Y(_00292_)
  );
  NAND3X1 _06665_ (
    .A(_00507_),
    .B(_00520_),
    .C(_00521_),
    .Y(_00524_)
  );
  NOR3X1 _06666_ (
    .A(_00513_),
    .B(_00516_),
    .C(_00524_),
    .Y(_00525_)
  );
  OAI21X1 _06667_ (
    .A(_00378_),
    .B(_00380_),
    .C(_00407_),
    .Y(_00526_)
  );
  INVX1 _06668_ (
    .A(_00526_),
    .Y(_00527_)
  );
  NOR2X1 _06669_ (
    .A(_00525_),
    .B(_00527_),
    .Y(_00528_)
  );
  XNOR2X1 _06670_ (
    .A(dbg_0.mem_cnt_8_ ),
    .B(_00407_),
    .Y(_00529_)
  );
  INVX1 _06671_ (
    .A(_00529_),
    .Y(_00530_)
  );
  OAI21X1 _06672_ (
    .A(_00525_),
    .B(_00527_),
    .C(_00530_),
    .Y(_00531_)
  );
  AOI21X1 _06673_ (
    .A(_00528_),
    .B(_00529_),
    .C(_00490_),
    .Y(_00532_)
  );
  OAI21X1 _06674_ (
    .A(_00528_),
    .B(_00529_),
    .C(_00532_),
    .Y(_00533_)
  );
  OAI21X1 _06675_ (
    .A(_00353_),
    .B(_00491_),
    .C(_00533_),
    .Y(_00293_)
  );
  NOR2X1 _06676_ (
    .A(dbg_0.dbg_din_9_ ),
    .B(_00491_),
    .Y(_00534_)
  );
  OAI21X1 _06677_ (
    .A(_00324_),
    .B(_00408_),
    .C(_00531_),
    .Y(_00535_)
  );
  XNOR2X1 _06678_ (
    .A(dbg_0.mem_cnt_9_ ),
    .B(_00407_),
    .Y(_00536_)
  );
  XOR2X1 _06679_ (
    .A(_00535_),
    .B(_00536_),
    .Y(_00537_)
  );
  AOI21X1 _06680_ (
    .A(_00491_),
    .B(_00537_),
    .C(_00534_),
    .Y(_00294_)
  );
  NAND2X1 _06681_ (
    .A(dbg_0.dbg_din_10_ ),
    .B(_00490_),
    .Y(_00538_)
  );
  OAI22X1 _06682_ (
    .A(_00373_),
    .B(_00408_),
    .C(_00531_),
    .D(_00536_),
    .Y(_00539_)
  );
  XNOR2X1 _06683_ (
    .A(dbg_0.mem_cnt_10_ ),
    .B(_00408_),
    .Y(_00540_)
  );
  AND2X1 _06684_ (
    .A(_00539_),
    .B(_00540_),
    .Y(_00541_)
  );
  OAI21X1 _06685_ (
    .A(_00539_),
    .B(_00540_),
    .C(_00491_),
    .Y(_00542_)
  );
  OAI21X1 _06686_ (
    .A(_00541_),
    .B(_00542_),
    .C(_00538_),
    .Y(_00280_)
  );
  AOI21X1 _06687_ (
    .A(dbg_0.mem_cnt_10_ ),
    .B(_00407_),
    .C(_00541_),
    .Y(_00543_)
  );
  XNOR2X1 _06688_ (
    .A(dbg_0.mem_cnt_11_ ),
    .B(_00408_),
    .Y(_00544_)
  );
  XOR2X1 _06689_ (
    .A(_00543_),
    .B(_00544_),
    .Y(_00545_)
  );
  MUX2X1 _06690_ (
    .A(_00357_),
    .B(_00545_),
    .S(_00490_),
    .Y(_00281_)
  );
  OAI21X1 _06691_ (
    .A(_00374_),
    .B(_00376_),
    .C(_00407_),
    .Y(_00546_)
  );
  INVX1 _06692_ (
    .A(_00546_),
    .Y(_00547_)
  );
  NAND2X1 _06693_ (
    .A(_00540_),
    .B(_00544_),
    .Y(_00548_)
  );
  NOR3X1 _06694_ (
    .A(_00531_),
    .B(_00536_),
    .C(_00548_),
    .Y(_00549_)
  );
  NOR2X1 _06695_ (
    .A(_00547_),
    .B(_00549_),
    .Y(_00550_)
  );
  OR2X1 _06696_ (
    .A(_00547_),
    .B(_00549_),
    .Y(_00551_)
  );
  XNOR2X1 _06697_ (
    .A(dbg_0.mem_cnt_12_ ),
    .B(_00407_),
    .Y(_00552_)
  );
  INVX1 _06698_ (
    .A(_00552_),
    .Y(_00553_)
  );
  AOI21X1 _06699_ (
    .A(_00550_),
    .B(_00552_),
    .C(_00490_),
    .Y(_00554_)
  );
  OAI21X1 _06700_ (
    .A(_00550_),
    .B(_00552_),
    .C(_00554_),
    .Y(_00555_)
  );
  OAI21X1 _06701_ (
    .A(_00359_),
    .B(_00491_),
    .C(_00555_),
    .Y(_00282_)
  );
  NOR2X1 _06702_ (
    .A(dbg_0.dbg_din_13_ ),
    .B(_00491_),
    .Y(_00556_)
  );
  AOI22X1 _06703_ (
    .A(dbg_0.mem_cnt_12_ ),
    .B(_00405_),
    .C(_00551_),
    .D(_00553_),
    .Y(_00557_)
  );
  NAND2X1 _06704_ (
    .A(dbg_0.mem_cnt_13_ ),
    .B(_00407_),
    .Y(_00558_)
  );
  XNOR2X1 _06705_ (
    .A(dbg_0.mem_cnt_13_ ),
    .B(_00407_),
    .Y(_00559_)
  );
  AND2X1 _06706_ (
    .A(_00557_),
    .B(_00558_),
    .Y(_00560_)
  );
  XNOR2X1 _06707_ (
    .A(_00557_),
    .B(_00559_),
    .Y(_00561_)
  );
  AOI21X1 _06708_ (
    .A(_00491_),
    .B(_00561_),
    .C(_00556_),
    .Y(_00283_)
  );
  NAND2X1 _06709_ (
    .A(dbg_0.mem_cnt_14_ ),
    .B(_00407_),
    .Y(_00562_)
  );
  XNOR2X1 _06710_ (
    .A(dbg_0.mem_cnt_14_ ),
    .B(_00407_),
    .Y(_00563_)
  );
  AOI21X1 _06711_ (
    .A(_00560_),
    .B(_00563_),
    .C(_00490_),
    .Y(_00564_)
  );
  OAI21X1 _06712_ (
    .A(_00560_),
    .B(_00563_),
    .C(_00564_),
    .Y(_00565_)
  );
  OAI21X1 _06713_ (
    .A(_00360_),
    .B(_00491_),
    .C(_00565_),
    .Y(_00284_)
  );
  OAI21X1 _06714_ (
    .A(_00560_),
    .B(_00563_),
    .C(_00562_),
    .Y(_00566_)
  );
  XNOR2X1 _06715_ (
    .A(dbg_0.mem_cnt_15_ ),
    .B(_00408_),
    .Y(_00567_)
  );
  XNOR2X1 _06716_ (
    .A(_00566_),
    .B(_00567_),
    .Y(_00568_)
  );
  NAND2X1 _06717_ (
    .A(dbg_0.dbg_din_15_ ),
    .B(_00490_),
    .Y(_00569_)
  );
  OAI21X1 _06718_ (
    .A(_00490_),
    .B(_00568_),
    .C(_00569_),
    .Y(_00285_)
  );
  NAND2X1 _06719_ (
    .A(dbg_0.dbg_din_0_ ),
    .B(_00486_),
    .Y(_00570_)
  );
  AND2X1 _06720_ (
    .A(dbg_en),
    .B(dbg_0.cpu_ctl_5_ ),
    .Y(_00571_)
  );
  AOI21X1 _06721_ (
    .A(_00162_),
    .B(_00571_),
    .C(dbg_0.halt_flag ),
    .Y(_00572_)
  );
  NAND2X1 _06722_ (
    .A(dbg_0.fe_mdb_in_1_ ),
    .B(dbg_0.fe_mdb_in_0_ ),
    .Y(_00573_)
  );
  NOR2X1 _06723_ (
    .A(dbg_0.fe_mdb_in_3_ ),
    .B(dbg_0.fe_mdb_in_2_ ),
    .Y(_00574_)
  );
  NOR2X1 _06724_ (
    .A(dbg_0.fe_mdb_in_5_ ),
    .B(dbg_0.fe_mdb_in_4_ ),
    .Y(_00575_)
  );
  NAND2X1 _06725_ (
    .A(_00574_),
    .B(_00575_),
    .Y(_00576_)
  );
  NOR2X1 _06726_ (
    .A(_00573_),
    .B(_00576_),
    .Y(_00577_)
  );
  NAND2X1 _06727_ (
    .A(_00363_),
    .B(dbg_0.fe_mdb_in_14_ ),
    .Y(_00578_)
  );
  NAND2X1 _06728_ (
    .A(dbg_0.decode_noirq ),
    .B(dbg_0.cpu_ctl_3_ ),
    .Y(_00579_)
  );
  NOR2X1 _06729_ (
    .A(_00578_),
    .B(_00579_),
    .Y(_00580_)
  );
  NOR2X1 _06730_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(dbg_0.fe_mdb_in_12_ ),
    .Y(_00581_)
  );
  NOR2X1 _06731_ (
    .A(dbg_0.fe_mdb_in_11_ ),
    .B(dbg_0.fe_mdb_in_10_ ),
    .Y(_00582_)
  );
  NAND2X1 _06732_ (
    .A(_00581_),
    .B(_00582_),
    .Y(_00583_)
  );
  NOR2X1 _06733_ (
    .A(dbg_0.fe_mdb_in_7_ ),
    .B(_00362_),
    .Y(_00584_)
  );
  NAND3X1 _06734_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(dbg_0.fe_mdb_in_8_ ),
    .C(_00584_),
    .Y(_00585_)
  );
  NOR2X1 _06735_ (
    .A(_00583_),
    .B(_00585_),
    .Y(_00586_)
  );
  NAND3X1 _06736_ (
    .A(_00577_),
    .B(_00580_),
    .C(_00586_),
    .Y(_00587_)
  );
  AND2X1 _06737_ (
    .A(_00572_),
    .B(_00587_),
    .Y(_00588_)
  );
  OAI21X1 _06738_ (
    .A(cpu_halt_st),
    .B(_00570_),
    .C(_00588_),
    .Y(_00589_)
  );
  AOI21X1 _06739_ (
    .A(dbg_0.mem_state_0_ ),
    .B(_00319_),
    .C(_00589_),
    .Y(_00590_)
  );
  NAND3X1 _06740_ (
    .A(cpu_halt_st),
    .B(dbg_0.dbg_din_1_ ),
    .C(_00486_),
    .Y(_00591_)
  );
  AOI21X1 _06741_ (
    .A(dbg_0.mem_state_1_ ),
    .B(_00395_),
    .C(_00590_),
    .Y(_00592_)
  );
  AND2X1 _06742_ (
    .A(_00591_),
    .B(_00592_),
    .Y(_00260_)
  );
  NAND2X1 _06743_ (
    .A(_00340_),
    .B(_00413_),
    .Y(_00593_)
  );
  NOR2X1 _06744_ (
    .A(_00417_),
    .B(_00593_),
    .Y(_00594_)
  );
  NOR2X1 _06745_ (
    .A(_00421_),
    .B(_00593_),
    .Y(_00595_)
  );
  NAND2X1 _06746_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00595_),
    .Y(_00596_)
  );
  NAND2X1 _06747_ (
    .A(_00328_),
    .B(_00596_),
    .Y(_00597_)
  );
  OAI21X1 _06748_ (
    .A(dbg_0.dbg_din_1_ ),
    .B(_00596_),
    .C(_00597_),
    .Y(_00598_)
  );
  INVX1 _06749_ (
    .A(_00598_),
    .Y(_00295_)
  );
  MUX2X1 _06750_ (
    .A(dbg_0.mem_ctl_2_ ),
    .B(dbg_0.dbg_din_2_ ),
    .S(_00596_),
    .Y(_00599_)
  );
  INVX1 _06751_ (
    .A(_00599_),
    .Y(_00296_)
  );
  MUX2X1 _06752_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(dbg_0.dbg_din_3_ ),
    .S(_00596_),
    .Y(_00600_)
  );
  INVX1 _06753_ (
    .A(_00600_),
    .Y(_00297_)
  );
  MUX2X1 _06754_ (
    .A(dbg_0.dbg_din_3_ ),
    .B(dbg_0.cpu_ctl_3_ ),
    .S(_00486_),
    .Y(_00601_)
  );
  INVX1 _06755_ (
    .A(_00601_),
    .Y(_00253_)
  );
  MUX2X1 _06756_ (
    .A(dbg_0.dbg_din_4_ ),
    .B(dbg_0.cpu_ctl_4_ ),
    .S(_00486_),
    .Y(_00602_)
  );
  INVX1 _06757_ (
    .A(_00602_),
    .Y(_00254_)
  );
  MUX2X1 _06758_ (
    .A(dbg_0.dbg_din_5_ ),
    .B(dbg_0.cpu_ctl_5_ ),
    .S(_00486_),
    .Y(_00603_)
  );
  INVX1 _06759_ (
    .A(_00603_),
    .Y(_00255_)
  );
  MUX2X1 _06760_ (
    .A(dbg_0.dbg_din_6_ ),
    .B(clock_module_0.dbg_cpu_reset ),
    .S(_00486_),
    .Y(_00604_)
  );
  INVX1 _06761_ (
    .A(_00604_),
    .Y(_00256_)
  );
  NOR2X1 _06762_ (
    .A(_00421_),
    .B(_00483_),
    .Y(_00605_)
  );
  AND2X1 _06763_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00605_),
    .Y(_00606_)
  );
  NAND2X1 _06764_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00605_),
    .Y(_00607_)
  );
  OAI21X1 _06765_ (
    .A(dbg_0.mem_ctl_1_ ),
    .B(_00479_),
    .C(dbg_0.dbg_mem_rd_dly ),
    .Y(_00608_)
  );
  MUX2X1 _06766_ (
    .A(dbg_0.dbg_mem_din_0_ ),
    .B(dbg_0.dbg_mem_din_8_ ),
    .S(_00393_),
    .Y(_00609_)
  );
  NAND2X1 _06767_ (
    .A(dbg_0.dbg_reg_din_0_ ),
    .B(_00480_),
    .Y(_00610_)
  );
  OAI21X1 _06768_ (
    .A(_00608_),
    .B(_00609_),
    .C(_00610_),
    .Y(_00611_)
  );
  AOI21X1 _06769_ (
    .A(dbg_0.mem_data_0_ ),
    .B(_00481_),
    .C(_00611_),
    .Y(_00612_)
  );
  NAND2X1 _06770_ (
    .A(dbg_0.dbg_din_0_ ),
    .B(_00606_),
    .Y(_00613_)
  );
  OAI21X1 _06771_ (
    .A(_00606_),
    .B(_00612_),
    .C(_00613_),
    .Y(_00298_)
  );
  MUX2X1 _06772_ (
    .A(dbg_0.dbg_mem_din_1_ ),
    .B(dbg_0.dbg_mem_din_9_ ),
    .S(_00393_),
    .Y(_00614_)
  );
  NAND2X1 _06773_ (
    .A(dbg_0.dbg_reg_din_1_ ),
    .B(_00480_),
    .Y(_00615_)
  );
  OAI21X1 _06774_ (
    .A(_00608_),
    .B(_00614_),
    .C(_00615_),
    .Y(_00616_)
  );
  AOI21X1 _06775_ (
    .A(dbg_0.mem_data_1_ ),
    .B(_00481_),
    .C(_00616_),
    .Y(_00617_)
  );
  NAND2X1 _06776_ (
    .A(dbg_0.dbg_din_1_ ),
    .B(_00606_),
    .Y(_00618_)
  );
  OAI21X1 _06777_ (
    .A(_00606_),
    .B(_00617_),
    .C(_00618_),
    .Y(_00305_)
  );
  NAND2X1 _06778_ (
    .A(dbg_0.mem_data_2_ ),
    .B(_00481_),
    .Y(_00619_)
  );
  AND2X1 _06779_ (
    .A(dbg_0.dbg_reg_din_2_ ),
    .B(_00480_),
    .Y(_00620_)
  );
  MUX2X1 _06780_ (
    .A(dbg_0.dbg_mem_din_2_ ),
    .B(dbg_0.dbg_mem_din_10_ ),
    .S(_00393_),
    .Y(_00621_)
  );
  OAI21X1 _06781_ (
    .A(_00608_),
    .B(_00621_),
    .C(_00619_),
    .Y(_00622_)
  );
  OAI21X1 _06782_ (
    .A(_00620_),
    .B(_00622_),
    .C(_00607_),
    .Y(_00623_)
  );
  OAI21X1 _06783_ (
    .A(_00343_),
    .B(_00607_),
    .C(_00623_),
    .Y(_00306_)
  );
  NAND2X1 _06784_ (
    .A(dbg_0.mem_data_3_ ),
    .B(_00481_),
    .Y(_00624_)
  );
  AND2X1 _06785_ (
    .A(dbg_0.dbg_reg_din_3_ ),
    .B(_00480_),
    .Y(_00625_)
  );
  MUX2X1 _06786_ (
    .A(dbg_0.dbg_mem_din_3_ ),
    .B(dbg_0.dbg_mem_din_11_ ),
    .S(_00393_),
    .Y(_00626_)
  );
  OAI21X1 _06787_ (
    .A(_00608_),
    .B(_00626_),
    .C(_00624_),
    .Y(_00627_)
  );
  OAI21X1 _06788_ (
    .A(_00625_),
    .B(_00627_),
    .C(_00607_),
    .Y(_00628_)
  );
  OAI21X1 _06789_ (
    .A(_00345_),
    .B(_00607_),
    .C(_00628_),
    .Y(_00307_)
  );
  NAND2X1 _06790_ (
    .A(dbg_0.dbg_reg_din_4_ ),
    .B(_00480_),
    .Y(_00629_)
  );
  MUX2X1 _06791_ (
    .A(dbg_0.dbg_mem_din_4_ ),
    .B(dbg_0.dbg_mem_din_12_ ),
    .S(_00393_),
    .Y(_00630_)
  );
  OAI21X1 _06792_ (
    .A(_00608_),
    .B(_00630_),
    .C(_00629_),
    .Y(_00631_)
  );
  AOI21X1 _06793_ (
    .A(dbg_0.mem_data_4_ ),
    .B(_00481_),
    .C(_00631_),
    .Y(_00632_)
  );
  NAND2X1 _06794_ (
    .A(dbg_0.dbg_din_4_ ),
    .B(_00606_),
    .Y(_00633_)
  );
  OAI21X1 _06795_ (
    .A(_00606_),
    .B(_00632_),
    .C(_00633_),
    .Y(_00308_)
  );
  NAND2X1 _06796_ (
    .A(dbg_0.dbg_reg_din_5_ ),
    .B(_00480_),
    .Y(_00634_)
  );
  MUX2X1 _06797_ (
    .A(dbg_0.dbg_mem_din_5_ ),
    .B(dbg_0.dbg_mem_din_13_ ),
    .S(_00393_),
    .Y(_00635_)
  );
  OAI21X1 _06798_ (
    .A(_00608_),
    .B(_00635_),
    .C(_00634_),
    .Y(_00636_)
  );
  AOI21X1 _06799_ (
    .A(dbg_0.mem_data_5_ ),
    .B(_00481_),
    .C(_00636_),
    .Y(_00637_)
  );
  NAND2X1 _06800_ (
    .A(dbg_0.dbg_din_5_ ),
    .B(_00606_),
    .Y(_00638_)
  );
  OAI21X1 _06801_ (
    .A(_00606_),
    .B(_00637_),
    .C(_00638_),
    .Y(_00309_)
  );
  NAND2X1 _06802_ (
    .A(dbg_0.dbg_reg_din_6_ ),
    .B(_00480_),
    .Y(_00639_)
  );
  MUX2X1 _06803_ (
    .A(dbg_0.dbg_mem_din_6_ ),
    .B(dbg_0.dbg_mem_din_14_ ),
    .S(_00393_),
    .Y(_00640_)
  );
  OAI21X1 _06804_ (
    .A(_00608_),
    .B(_00640_),
    .C(_00639_),
    .Y(_00641_)
  );
  AOI21X1 _06805_ (
    .A(dbg_0.mem_data_6_ ),
    .B(_00481_),
    .C(_00641_),
    .Y(_00642_)
  );
  NAND2X1 _06806_ (
    .A(dbg_0.dbg_din_6_ ),
    .B(_00606_),
    .Y(_00643_)
  );
  OAI21X1 _06807_ (
    .A(_00606_),
    .B(_00642_),
    .C(_00643_),
    .Y(_00310_)
  );
  NAND2X1 _06808_ (
    .A(dbg_0.mem_data_7_ ),
    .B(_00481_),
    .Y(_00644_)
  );
  MUX2X1 _06809_ (
    .A(dbg_0.dbg_mem_din_7_ ),
    .B(dbg_0.dbg_mem_din_15_ ),
    .S(_00393_),
    .Y(_00645_)
  );
  AND2X1 _06810_ (
    .A(dbg_0.dbg_reg_din_7_ ),
    .B(_00480_),
    .Y(_00646_)
  );
  OAI21X1 _06811_ (
    .A(_00608_),
    .B(_00645_),
    .C(_00644_),
    .Y(_00647_)
  );
  OAI21X1 _06812_ (
    .A(_00646_),
    .B(_00647_),
    .C(_00607_),
    .Y(_00648_)
  );
  OAI21X1 _06813_ (
    .A(_00351_),
    .B(_00607_),
    .C(_00648_),
    .Y(_00311_)
  );
  NOR2X1 _06814_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00361_),
    .Y(_00649_)
  );
  NAND2X1 _06815_ (
    .A(dbg_0.dbg_mem_din_8_ ),
    .B(_00649_),
    .Y(_00650_)
  );
  NAND2X1 _06816_ (
    .A(dbg_0.dbg_reg_din_8_ ),
    .B(_00480_),
    .Y(_00651_)
  );
  OAI21X1 _06817_ (
    .A(_00480_),
    .B(_00650_),
    .C(_00651_),
    .Y(_00652_)
  );
  AOI21X1 _06818_ (
    .A(dbg_0.mem_data_8_ ),
    .B(_00481_),
    .C(_00652_),
    .Y(_00653_)
  );
  MUX2X1 _06819_ (
    .A(_00353_),
    .B(_00653_),
    .S(_00606_),
    .Y(_00312_)
  );
  NAND2X1 _06820_ (
    .A(dbg_0.dbg_mem_din_9_ ),
    .B(_00649_),
    .Y(_00654_)
  );
  NAND2X1 _06821_ (
    .A(dbg_0.dbg_reg_din_9_ ),
    .B(_00480_),
    .Y(_00655_)
  );
  OAI21X1 _06822_ (
    .A(_00480_),
    .B(_00654_),
    .C(_00655_),
    .Y(_00656_)
  );
  AOI21X1 _06823_ (
    .A(dbg_0.mem_data_9_ ),
    .B(_00481_),
    .C(_00656_),
    .Y(_00657_)
  );
  NOR2X1 _06824_ (
    .A(dbg_0.dbg_din_9_ ),
    .B(_00607_),
    .Y(_00658_)
  );
  AOI21X1 _06825_ (
    .A(_00607_),
    .B(_00657_),
    .C(_00658_),
    .Y(_00313_)
  );
  NAND2X1 _06826_ (
    .A(dbg_0.dbg_mem_din_10_ ),
    .B(_00649_),
    .Y(_00659_)
  );
  NAND2X1 _06827_ (
    .A(dbg_0.dbg_reg_din_10_ ),
    .B(_00480_),
    .Y(_00660_)
  );
  OAI21X1 _06828_ (
    .A(_00480_),
    .B(_00659_),
    .C(_00660_),
    .Y(_00661_)
  );
  AOI21X1 _06829_ (
    .A(dbg_0.mem_data_10_ ),
    .B(_00481_),
    .C(_00661_),
    .Y(_00662_)
  );
  NOR2X1 _06830_ (
    .A(dbg_0.dbg_din_10_ ),
    .B(_00607_),
    .Y(_00663_)
  );
  AOI21X1 _06831_ (
    .A(_00607_),
    .B(_00662_),
    .C(_00663_),
    .Y(_00299_)
  );
  NAND2X1 _06832_ (
    .A(dbg_0.dbg_mem_din_11_ ),
    .B(_00649_),
    .Y(_00664_)
  );
  NAND2X1 _06833_ (
    .A(dbg_0.dbg_reg_din_11_ ),
    .B(_00480_),
    .Y(_00665_)
  );
  OAI21X1 _06834_ (
    .A(_00480_),
    .B(_00664_),
    .C(_00665_),
    .Y(_00666_)
  );
  AOI21X1 _06835_ (
    .A(dbg_0.mem_data_11_ ),
    .B(_00481_),
    .C(_00666_),
    .Y(_00667_)
  );
  MUX2X1 _06836_ (
    .A(_00357_),
    .B(_00667_),
    .S(_00606_),
    .Y(_00300_)
  );
  NAND2X1 _06837_ (
    .A(dbg_0.dbg_mem_din_12_ ),
    .B(_00649_),
    .Y(_00668_)
  );
  NAND2X1 _06838_ (
    .A(dbg_0.dbg_reg_din_12_ ),
    .B(_00480_),
    .Y(_00669_)
  );
  OAI21X1 _06839_ (
    .A(_00480_),
    .B(_00668_),
    .C(_00669_),
    .Y(_00670_)
  );
  AOI21X1 _06840_ (
    .A(dbg_0.mem_data_12_ ),
    .B(_00481_),
    .C(_00670_),
    .Y(_00671_)
  );
  MUX2X1 _06841_ (
    .A(_00359_),
    .B(_00671_),
    .S(_00606_),
    .Y(_00301_)
  );
  NAND2X1 _06842_ (
    .A(dbg_0.dbg_mem_din_13_ ),
    .B(_00649_),
    .Y(_00672_)
  );
  NAND2X1 _06843_ (
    .A(dbg_0.dbg_reg_din_13_ ),
    .B(_00480_),
    .Y(_00673_)
  );
  OAI21X1 _06844_ (
    .A(_00480_),
    .B(_00672_),
    .C(_00673_),
    .Y(_00674_)
  );
  AOI21X1 _06845_ (
    .A(dbg_0.mem_data_13_ ),
    .B(_00481_),
    .C(_00674_),
    .Y(_00675_)
  );
  NOR2X1 _06846_ (
    .A(dbg_0.dbg_din_13_ ),
    .B(_00607_),
    .Y(_00676_)
  );
  AOI21X1 _06847_ (
    .A(_00607_),
    .B(_00675_),
    .C(_00676_),
    .Y(_00302_)
  );
  NAND2X1 _06848_ (
    .A(dbg_0.dbg_mem_din_14_ ),
    .B(_00649_),
    .Y(_00677_)
  );
  NAND2X1 _06849_ (
    .A(dbg_0.dbg_reg_din_14_ ),
    .B(_00480_),
    .Y(_00678_)
  );
  OAI21X1 _06850_ (
    .A(_00480_),
    .B(_00677_),
    .C(_00678_),
    .Y(_00679_)
  );
  AOI21X1 _06851_ (
    .A(dbg_0.mem_data_14_ ),
    .B(_00481_),
    .C(_00679_),
    .Y(_00680_)
  );
  MUX2X1 _06852_ (
    .A(_00360_),
    .B(_00680_),
    .S(_00606_),
    .Y(_00303_)
  );
  NAND2X1 _06853_ (
    .A(dbg_0.dbg_mem_din_15_ ),
    .B(_00649_),
    .Y(_00681_)
  );
  NAND2X1 _06854_ (
    .A(dbg_0.dbg_reg_din_15_ ),
    .B(_00480_),
    .Y(_00682_)
  );
  OAI21X1 _06855_ (
    .A(_00480_),
    .B(_00681_),
    .C(_00682_),
    .Y(_00683_)
  );
  AOI21X1 _06856_ (
    .A(dbg_0.mem_data_15_ ),
    .B(_00481_),
    .C(_00683_),
    .Y(_00684_)
  );
  NOR2X1 _06857_ (
    .A(dbg_0.dbg_din_15_ ),
    .B(_00607_),
    .Y(_00685_)
  );
  AOI21X1 _06858_ (
    .A(_00607_),
    .B(_00684_),
    .C(_00685_),
    .Y(_00304_)
  );
  NOR2X1 _06859_ (
    .A(_00484_),
    .B(_00488_),
    .Y(_00686_)
  );
  NAND2X1 _06860_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00686_),
    .Y(_00687_)
  );
  OR2X1 _06861_ (
    .A(_00343_),
    .B(_00687_),
    .Y(_00688_)
  );
  AOI21X1 _06862_ (
    .A(dbg_0.cpu_stat_2_ ),
    .B(_00688_),
    .C(_00162_),
    .Y(_00689_)
  );
  INVX1 _06863_ (
    .A(_00689_),
    .Y(_00257_)
  );
  OAI21X1 _06864_ (
    .A(_00345_),
    .B(_00687_),
    .C(dbg_0.cpu_stat_3_ ),
    .Y(_00690_)
  );
  NAND2X1 _06865_ (
    .A(_00587_),
    .B(_00690_),
    .Y(_00258_)
  );
  NAND3X1 _06866_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(dbg_0.dbg_din_0_ ),
    .C(_00594_),
    .Y(_00691_)
  );
  INVX1 _06867_ (
    .A(_00691_),
    .Y(_00314_)
  );
  NOR2X1 _06868_ (
    .A(_00328_),
    .B(_00479_),
    .Y(dbg_0.dbg_reg_wr )
  );
  NOR2X1 _06869_ (
    .A(_00414_),
    .B(_00484_),
    .Y(_00692_)
  );
  NOR2X1 _06870_ (
    .A(_00484_),
    .B(_00593_),
    .Y(_00693_)
  );
  NAND2X1 _06871_ (
    .A(dbg_0.dbg_addr_3_ ),
    .B(dbg_0.dbg_addr_4_ ),
    .Y(_00694_)
  );
  NOR2X1 _06872_ (
    .A(dbg_0.dbg_addr_5_ ),
    .B(_00694_),
    .Y(_00695_)
  );
  NAND2X1 _06873_ (
    .A(_00420_),
    .B(_00695_),
    .Y(_00696_)
  );
  NOR2X1 _06874_ (
    .A(_00593_),
    .B(_00696_),
    .Y(_00697_)
  );
  AOI22X1 _06875_ (
    .A(cpu_halt_st),
    .B(_00686_),
    .C(_00692_),
    .D(1'h1),
    .Y(_00698_)
  );
  INVX1 _06876_ (
    .A(_00698_),
    .Y(_00699_)
  );
  AOI21X1 _06877_ (
    .A(dbg_0.mem_data_0_ ),
    .B(_00605_),
    .C(_00699_),
    .Y(_00700_)
  );
  AOI22X1 _06878_ (
    .A(dbg_0.dbg_mem_addr_0_ ),
    .B(_00422_),
    .C(_00697_),
    .D(1'h0),
    .Y(_00701_)
  );
  AOI22X1 _06879_ (
    .A(dbg_0.mem_cnt_0_ ),
    .B(_00489_),
    .C(_00693_),
    .D(1'h1),
    .Y(_00702_)
  );
  NAND3X1 _06880_ (
    .A(_00700_),
    .B(_00701_),
    .C(_00702_),
    .Y(dbg_0.dbg_dout_0_ )
  );
  AOI22X1 _06881_ (
    .A(dbg_0.dbg_mem_addr_1_ ),
    .B(_00422_),
    .C(_00693_),
    .D(1'h1),
    .Y(_00703_)
  );
  AOI22X1 _06882_ (
    .A(dbg_0.mem_cnt_1_ ),
    .B(_00489_),
    .C(_00692_),
    .D(1'h0),
    .Y(_00704_)
  );
  AOI22X1 _06883_ (
    .A(dbg_0.mem_ctl_1_ ),
    .B(_00595_),
    .C(_00697_),
    .D(1'h0),
    .Y(_00705_)
  );
  INVX1 _06884_ (
    .A(_00705_),
    .Y(_00706_)
  );
  AOI21X1 _06885_ (
    .A(dbg_0.mem_data_1_ ),
    .B(_00605_),
    .C(_00706_),
    .Y(_00707_)
  );
  NAND3X1 _06886_ (
    .A(_00703_),
    .B(_00704_),
    .C(_00707_),
    .Y(dbg_0.dbg_dout_1_ )
  );
  NAND2X1 _06887_ (
    .A(dbg_0.cpu_stat_2_ ),
    .B(_00686_),
    .Y(_00708_)
  );
  AOI22X1 _06888_ (
    .A(dbg_0.dbg_mem_addr_2_ ),
    .B(_00418_),
    .C(_00594_),
    .D(dbg_0.mem_ctl_2_ ),
    .Y(_00709_)
  );
  AOI22X1 _06889_ (
    .A(1'h0),
    .B(_00693_),
    .C(_00697_),
    .D(1'h0),
    .Y(_00710_)
  );
  AOI22X1 _06890_ (
    .A(dbg_0.mem_cnt_2_ ),
    .B(_00489_),
    .C(_00692_),
    .D(1'h0),
    .Y(_00711_)
  );
  NAND2X1 _06891_ (
    .A(_00710_),
    .B(_00711_),
    .Y(_00712_)
  );
  AOI21X1 _06892_ (
    .A(dbg_0.mem_data_2_ ),
    .B(_00605_),
    .C(_00712_),
    .Y(_00713_)
  );
  NAND3X1 _06893_ (
    .A(_00708_),
    .B(_00709_),
    .C(_00713_),
    .Y(dbg_0.dbg_dout_2_ )
  );
  AOI22X1 _06894_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00595_),
    .C(_00697_),
    .D(1'h0),
    .Y(_00714_)
  );
  AOI22X1 _06895_ (
    .A(dbg_0.cpu_ctl_3_ ),
    .B(_00485_),
    .C(_00692_),
    .D(1'h0),
    .Y(_00715_)
  );
  AOI22X1 _06896_ (
    .A(dbg_0.mem_cnt_3_ ),
    .B(_00489_),
    .C(_00693_),
    .D(1'h0),
    .Y(_00716_)
  );
  AOI22X1 _06897_ (
    .A(dbg_0.dbg_mem_addr_3_ ),
    .B(_00418_),
    .C(_00686_),
    .D(dbg_0.cpu_stat_3_ ),
    .Y(_00717_)
  );
  NAND2X1 _06898_ (
    .A(_00716_),
    .B(_00717_),
    .Y(_00718_)
  );
  AOI21X1 _06899_ (
    .A(dbg_0.mem_data_3_ ),
    .B(_00605_),
    .C(_00718_),
    .Y(_00719_)
  );
  NAND3X1 _06900_ (
    .A(_00714_),
    .B(_00715_),
    .C(_00719_),
    .Y(dbg_0.dbg_dout_3_ )
  );
  AOI22X1 _06901_ (
    .A(dbg_0.cpu_ctl_4_ ),
    .B(_00485_),
    .C(_00489_),
    .D(dbg_0.mem_cnt_4_ ),
    .Y(_00720_)
  );
  AOI22X1 _06902_ (
    .A(1'h0),
    .B(_00692_),
    .C(_00693_),
    .D(1'h0),
    .Y(_00721_)
  );
  AOI22X1 _06903_ (
    .A(dbg_0.mem_data_4_ ),
    .B(_00605_),
    .C(_00697_),
    .D(1'h0),
    .Y(_00722_)
  );
  INVX1 _06904_ (
    .A(_00722_),
    .Y(_00723_)
  );
  AOI21X1 _06905_ (
    .A(dbg_0.dbg_mem_addr_4_ ),
    .B(_00422_),
    .C(_00723_),
    .Y(_00724_)
  );
  NAND3X1 _06906_ (
    .A(_00720_),
    .B(_00721_),
    .C(_00724_),
    .Y(dbg_0.dbg_dout_4_ )
  );
  AOI22X1 _06907_ (
    .A(1'h0),
    .B(_00693_),
    .C(_00697_),
    .D(1'h0),
    .Y(_00725_)
  );
  AOI22X1 _06908_ (
    .A(dbg_0.mem_cnt_5_ ),
    .B(_00489_),
    .C(_00605_),
    .D(dbg_0.mem_data_5_ ),
    .Y(_00726_)
  );
  INVX1 _06909_ (
    .A(_00726_),
    .Y(_00727_)
  );
  AOI21X1 _06910_ (
    .A(dbg_0.cpu_ctl_5_ ),
    .B(_00485_),
    .C(_00727_),
    .Y(_00728_)
  );
  AOI22X1 _06911_ (
    .A(dbg_0.dbg_mem_addr_5_ ),
    .B(_00422_),
    .C(_00692_),
    .D(1'h0),
    .Y(_00729_)
  );
  NAND3X1 _06912_ (
    .A(_00725_),
    .B(_00728_),
    .C(_00729_),
    .Y(dbg_0.dbg_dout_5_ )
  );
  AOI22X1 _06913_ (
    .A(dbg_0.dbg_mem_addr_6_ ),
    .B(_00422_),
    .C(_00697_),
    .D(1'h0),
    .Y(_00730_)
  );
  INVX1 _06914_ (
    .A(_00730_),
    .Y(_00731_)
  );
  AOI21X1 _06915_ (
    .A(1'h0),
    .B(_00693_),
    .C(_00731_),
    .Y(_00732_)
  );
  AOI22X1 _06916_ (
    .A(clock_module_0.dbg_cpu_reset ),
    .B(_00485_),
    .C(_00692_),
    .D(1'h0),
    .Y(_00733_)
  );
  AOI22X1 _06917_ (
    .A(dbg_0.mem_cnt_6_ ),
    .B(_00489_),
    .C(_00605_),
    .D(dbg_0.mem_data_6_ ),
    .Y(_00734_)
  );
  NAND3X1 _06918_ (
    .A(_00732_),
    .B(_00733_),
    .C(_00734_),
    .Y(dbg_0.dbg_dout_6_ )
  );
  NAND2X1 _06919_ (
    .A(1'h0),
    .B(_00697_),
    .Y(_00735_)
  );
  AOI22X1 _06920_ (
    .A(dbg_0.dbg_mem_addr_7_ ),
    .B(_00422_),
    .C(_00692_),
    .D(1'h0),
    .Y(_00736_)
  );
  AOI22X1 _06921_ (
    .A(dbg_0.mem_cnt_7_ ),
    .B(_00489_),
    .C(_00605_),
    .D(dbg_0.mem_data_7_ ),
    .Y(_00737_)
  );
  INVX1 _06922_ (
    .A(_00737_),
    .Y(_00738_)
  );
  AOI21X1 _06923_ (
    .A(1'h0),
    .B(_00693_),
    .C(_00738_),
    .Y(_00739_)
  );
  NAND3X1 _06924_ (
    .A(_00735_),
    .B(_00736_),
    .C(_00739_),
    .Y(dbg_0.dbg_dout_7_ )
  );
  NAND2X1 _06925_ (
    .A(1'h0),
    .B(_00697_),
    .Y(_00740_)
  );
  AOI22X1 _06926_ (
    .A(dbg_0.mem_cnt_8_ ),
    .B(_00489_),
    .C(_00605_),
    .D(dbg_0.mem_data_8_ ),
    .Y(_00741_)
  );
  INVX1 _06927_ (
    .A(_00741_),
    .Y(_00742_)
  );
  AOI21X1 _06928_ (
    .A(1'h0),
    .B(_00693_),
    .C(_00742_),
    .Y(_00743_)
  );
  AOI22X1 _06929_ (
    .A(dbg_0.dbg_mem_addr_8_ ),
    .B(_00422_),
    .C(_00692_),
    .D(1'h1),
    .Y(_00744_)
  );
  NAND3X1 _06930_ (
    .A(_00740_),
    .B(_00743_),
    .C(_00744_),
    .Y(dbg_0.dbg_dout_8_ )
  );
  NAND2X1 _06931_ (
    .A(1'h0),
    .B(_00697_),
    .Y(_00745_)
  );
  AOI22X1 _06932_ (
    .A(dbg_0.mem_cnt_9_ ),
    .B(_00489_),
    .C(_00605_),
    .D(dbg_0.mem_data_9_ ),
    .Y(_00746_)
  );
  AOI22X1 _06933_ (
    .A(dbg_0.dbg_mem_addr_9_ ),
    .B(_00422_),
    .C(_00692_),
    .D(1'h0),
    .Y(_00747_)
  );
  INVX1 _06934_ (
    .A(_00747_),
    .Y(_00748_)
  );
  AOI21X1 _06935_ (
    .A(1'h0),
    .B(_00693_),
    .C(_00748_),
    .Y(_00749_)
  );
  NAND3X1 _06936_ (
    .A(_00745_),
    .B(_00746_),
    .C(_00749_),
    .Y(dbg_0.dbg_dout_9_ )
  );
  NAND2X1 _06937_ (
    .A(1'h0),
    .B(_00697_),
    .Y(_00750_)
  );
  AOI22X1 _06938_ (
    .A(dbg_0.dbg_mem_addr_10_ ),
    .B(_00422_),
    .C(_00489_),
    .D(dbg_0.mem_cnt_10_ ),
    .Y(_00751_)
  );
  AOI22X1 _06939_ (
    .A(1'h0),
    .B(_00692_),
    .C(_00693_),
    .D(1'h0),
    .Y(_00752_)
  );
  INVX1 _06940_ (
    .A(_00752_),
    .Y(_00753_)
  );
  AOI21X1 _06941_ (
    .A(dbg_0.mem_data_10_ ),
    .B(_00605_),
    .C(_00753_),
    .Y(_00754_)
  );
  NAND3X1 _06942_ (
    .A(_00750_),
    .B(_00751_),
    .C(_00754_),
    .Y(dbg_0.dbg_dout_10_ )
  );
  AOI22X1 _06943_ (
    .A(dbg_0.dbg_mem_addr_11_ ),
    .B(_00422_),
    .C(_00692_),
    .D(1'h0),
    .Y(_00755_)
  );
  INVX1 _06944_ (
    .A(_00755_),
    .Y(_00756_)
  );
  AOI21X1 _06945_ (
    .A(1'h0),
    .B(_00693_),
    .C(_00756_),
    .Y(_00757_)
  );
  NAND2X1 _06946_ (
    .A(dbg_0.mem_data_11_ ),
    .B(_00605_),
    .Y(_00758_)
  );
  AOI22X1 _06947_ (
    .A(dbg_0.mem_cnt_11_ ),
    .B(_00489_),
    .C(_00697_),
    .D(1'h0),
    .Y(_00759_)
  );
  NAND3X1 _06948_ (
    .A(_00757_),
    .B(_00758_),
    .C(_00759_),
    .Y(dbg_0.dbg_dout_11_ )
  );
  NAND2X1 _06949_ (
    .A(1'h0),
    .B(_00697_),
    .Y(_00760_)
  );
  AOI22X1 _06950_ (
    .A(dbg_0.mem_cnt_12_ ),
    .B(_00489_),
    .C(_00605_),
    .D(dbg_0.mem_data_12_ ),
    .Y(_00761_)
  );
  AOI22X1 _06951_ (
    .A(dbg_0.dbg_mem_addr_12_ ),
    .B(_00422_),
    .C(_00692_),
    .D(1'h0),
    .Y(_00762_)
  );
  INVX1 _06952_ (
    .A(_00762_),
    .Y(_00763_)
  );
  AOI21X1 _06953_ (
    .A(1'h0),
    .B(_00693_),
    .C(_00763_),
    .Y(_00764_)
  );
  NAND3X1 _06954_ (
    .A(_00760_),
    .B(_00761_),
    .C(_00764_),
    .Y(dbg_0.dbg_dout_12_ )
  );
  NAND2X1 _06955_ (
    .A(1'h0),
    .B(_00697_),
    .Y(_00765_)
  );
  AOI22X1 _06956_ (
    .A(dbg_0.mem_cnt_13_ ),
    .B(_00489_),
    .C(_00605_),
    .D(dbg_0.mem_data_13_ ),
    .Y(_00766_)
  );
  AOI22X1 _06957_ (
    .A(dbg_0.dbg_mem_addr_13_ ),
    .B(_00422_),
    .C(_00692_),
    .D(1'h0),
    .Y(_00767_)
  );
  INVX1 _06958_ (
    .A(_00767_),
    .Y(_00768_)
  );
  AOI21X1 _06959_ (
    .A(1'h0),
    .B(_00693_),
    .C(_00768_),
    .Y(_00769_)
  );
  NAND3X1 _06960_ (
    .A(_00765_),
    .B(_00766_),
    .C(_00769_),
    .Y(dbg_0.dbg_dout_13_ )
  );
  NAND2X1 _06961_ (
    .A(1'h0),
    .B(_00697_),
    .Y(_00770_)
  );
  AOI22X1 _06962_ (
    .A(dbg_0.dbg_mem_addr_14_ ),
    .B(_00422_),
    .C(_00489_),
    .D(dbg_0.mem_cnt_14_ ),
    .Y(_00771_)
  );
  INVX1 _06963_ (
    .A(_00771_),
    .Y(_00772_)
  );
  AOI21X1 _06964_ (
    .A(dbg_0.mem_data_14_ ),
    .B(_00605_),
    .C(_00772_),
    .Y(_00773_)
  );
  AOI22X1 _06965_ (
    .A(1'h0),
    .B(_00692_),
    .C(_00693_),
    .D(1'h1),
    .Y(_00774_)
  );
  NAND3X1 _06966_ (
    .A(_00770_),
    .B(_00773_),
    .C(_00774_),
    .Y(dbg_0.dbg_dout_14_ )
  );
  NAND2X1 _06967_ (
    .A(1'h0),
    .B(_00697_),
    .Y(_00775_)
  );
  AOI22X1 _06968_ (
    .A(dbg_0.dbg_mem_addr_15_ ),
    .B(_00422_),
    .C(_00692_),
    .D(1'h1),
    .Y(_00776_)
  );
  AOI22X1 _06969_ (
    .A(dbg_0.mem_cnt_15_ ),
    .B(_00489_),
    .C(_00605_),
    .D(dbg_0.mem_data_15_ ),
    .Y(_00777_)
  );
  INVX1 _06970_ (
    .A(_00777_),
    .Y(_00778_)
  );
  AOI21X1 _06971_ (
    .A(1'h0),
    .B(_00693_),
    .C(_00778_),
    .Y(_00779_)
  );
  NAND3X1 _06972_ (
    .A(_00775_),
    .B(_00776_),
    .C(_00779_),
    .Y(dbg_0.dbg_dout_15_ )
  );
  OAI21X1 _06973_ (
    .A(dbg_0.cpu_ctl_4_ ),
    .B(_00364_),
    .C(cpu_halt_st),
    .Y(_00780_)
  );
  INVX1 _06974_ (
    .A(_00780_),
    .Y(_00049_)
  );
  NOR2X1 _06975_ (
    .A(dbg_0.inc_step_1_ ),
    .B(_00590_),
    .Y(cpu_halt_cmd)
  );
  NOR2X1 _06976_ (
    .A(_00328_),
    .B(_00477_),
    .Y(dbg_0.dbg_i2c_0.mem_burst_wr )
  );
  OAI21X1 _06977_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(dbg_0.dbg_i2c_0.dbg_rd ),
    .C(dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00781_)
  );
  OAI21X1 _06978_ (
    .A(dbg_0.mem_ctl_1_ ),
    .B(_00477_),
    .C(_00781_),
    .Y(_00315_)
  );
  AND2X1 _06979_ (
    .A(_00328_),
    .B(dbg_0.dbg_mem_en ),
    .Y(dbg_0.dbg_mem_rd )
  );
  AOI21X1 _06980_ (
    .A(_00339_),
    .B(_00477_),
    .C(dbg_0.dbg_i2c_0.mem_burst_end ),
    .Y(_00278_)
  );
  DFFSR _06981_ (
    .CLK(dco_clk),
    .D(_00318_),
    .Q(dbg_0.mem_state_0_ ),
    .R(1'h1),
    .S(_00320_)
  );
  DFFSR _06982_ (
    .CLK(dco_clk),
    .D(_00316_),
    .Q(dbg_0.mem_state_1_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06983_ (
    .CLK(dco_clk),
    .D(_00319_),
    .Q(dbg_0.mem_state_2_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06984_ (
    .CLK(dco_clk),
    .D(_00317_),
    .Q(dbg_0.mem_state_3_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06985_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_mem_rd ),
    .Q(dbg_0.dbg_mem_rd_dly ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06986_ (
    .CLK(dco_clk),
    .D(_00315_),
    .Q(dbg_0.mem_startb ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06987_ (
    .CLK(dco_clk),
    .D(_00278_),
    .Q(dbg_0.dbg_i2c_0.mem_burst ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06988_ (
    .CLK(dco_clk),
    .D(_00260_),
    .Q(dbg_0.halt_flag ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06989_ (
    .CLK(dco_clk),
    .D(dbg_0.istep ),
    .Q(dbg_0.inc_step_0_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06990_ (
    .CLK(dco_clk),
    .D(_00261_),
    .Q(dbg_0.inc_step_1_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06991_ (
    .CLK(dco_clk),
    .D(_00259_),
    .Q(dbg_0.dbg_rd_rdy ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06992_ (
    .CLK(dco_clk),
    .D(_00279_),
    .Q(dbg_0.mem_cnt_0_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06993_ (
    .CLK(dco_clk),
    .D(_00286_),
    .Q(dbg_0.mem_cnt_1_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06994_ (
    .CLK(dco_clk),
    .D(_00287_),
    .Q(dbg_0.mem_cnt_2_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06995_ (
    .CLK(dco_clk),
    .D(_00288_),
    .Q(dbg_0.mem_cnt_3_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06996_ (
    .CLK(dco_clk),
    .D(_00289_),
    .Q(dbg_0.mem_cnt_4_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06997_ (
    .CLK(dco_clk),
    .D(_00290_),
    .Q(dbg_0.mem_cnt_5_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06998_ (
    .CLK(dco_clk),
    .D(_00291_),
    .Q(dbg_0.mem_cnt_6_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06999_ (
    .CLK(dco_clk),
    .D(_00292_),
    .Q(dbg_0.mem_cnt_7_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07000_ (
    .CLK(dco_clk),
    .D(_00293_),
    .Q(dbg_0.mem_cnt_8_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07001_ (
    .CLK(dco_clk),
    .D(_00294_),
    .Q(dbg_0.mem_cnt_9_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07002_ (
    .CLK(dco_clk),
    .D(_00280_),
    .Q(dbg_0.mem_cnt_10_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07003_ (
    .CLK(dco_clk),
    .D(_00281_),
    .Q(dbg_0.mem_cnt_11_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07004_ (
    .CLK(dco_clk),
    .D(_00282_),
    .Q(dbg_0.mem_cnt_12_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07005_ (
    .CLK(dco_clk),
    .D(_00283_),
    .Q(dbg_0.mem_cnt_13_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07006_ (
    .CLK(dco_clk),
    .D(_00284_),
    .Q(dbg_0.mem_cnt_14_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07007_ (
    .CLK(dco_clk),
    .D(_00285_),
    .Q(dbg_0.mem_cnt_15_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07008_ (
    .CLK(dco_clk),
    .D(_00262_),
    .Q(dbg_0.dbg_mem_addr_0_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07009_ (
    .CLK(dco_clk),
    .D(_00269_),
    .Q(dbg_0.dbg_mem_addr_1_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07010_ (
    .CLK(dco_clk),
    .D(_00270_),
    .Q(dbg_0.dbg_mem_addr_2_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07011_ (
    .CLK(dco_clk),
    .D(_00271_),
    .Q(dbg_0.dbg_mem_addr_3_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07012_ (
    .CLK(dco_clk),
    .D(_00272_),
    .Q(dbg_0.dbg_mem_addr_4_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07013_ (
    .CLK(dco_clk),
    .D(_00273_),
    .Q(dbg_0.dbg_mem_addr_5_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07014_ (
    .CLK(dco_clk),
    .D(_00274_),
    .Q(dbg_0.dbg_mem_addr_6_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07015_ (
    .CLK(dco_clk),
    .D(_00275_),
    .Q(dbg_0.dbg_mem_addr_7_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07016_ (
    .CLK(dco_clk),
    .D(_00276_),
    .Q(dbg_0.dbg_mem_addr_8_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07017_ (
    .CLK(dco_clk),
    .D(_00277_),
    .Q(dbg_0.dbg_mem_addr_9_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07018_ (
    .CLK(dco_clk),
    .D(_00263_),
    .Q(dbg_0.dbg_mem_addr_10_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07019_ (
    .CLK(dco_clk),
    .D(_00264_),
    .Q(dbg_0.dbg_mem_addr_11_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07020_ (
    .CLK(dco_clk),
    .D(_00265_),
    .Q(dbg_0.dbg_mem_addr_12_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07021_ (
    .CLK(dco_clk),
    .D(_00266_),
    .Q(dbg_0.dbg_mem_addr_13_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07022_ (
    .CLK(dco_clk),
    .D(_00267_),
    .Q(dbg_0.dbg_mem_addr_14_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07023_ (
    .CLK(dco_clk),
    .D(_00268_),
    .Q(dbg_0.dbg_mem_addr_15_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07024_ (
    .CLK(dco_clk),
    .D(_00298_),
    .Q(dbg_0.mem_data_0_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07025_ (
    .CLK(dco_clk),
    .D(_00305_),
    .Q(dbg_0.mem_data_1_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07026_ (
    .CLK(dco_clk),
    .D(_00306_),
    .Q(dbg_0.mem_data_2_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07027_ (
    .CLK(dco_clk),
    .D(_00307_),
    .Q(dbg_0.mem_data_3_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07028_ (
    .CLK(dco_clk),
    .D(_00308_),
    .Q(dbg_0.mem_data_4_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07029_ (
    .CLK(dco_clk),
    .D(_00309_),
    .Q(dbg_0.mem_data_5_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07030_ (
    .CLK(dco_clk),
    .D(_00310_),
    .Q(dbg_0.mem_data_6_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07031_ (
    .CLK(dco_clk),
    .D(_00311_),
    .Q(dbg_0.mem_data_7_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07032_ (
    .CLK(dco_clk),
    .D(_00312_),
    .Q(dbg_0.mem_data_8_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07033_ (
    .CLK(dco_clk),
    .D(_00313_),
    .Q(dbg_0.mem_data_9_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07034_ (
    .CLK(dco_clk),
    .D(_00299_),
    .Q(dbg_0.mem_data_10_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07035_ (
    .CLK(dco_clk),
    .D(_00300_),
    .Q(dbg_0.mem_data_11_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07036_ (
    .CLK(dco_clk),
    .D(_00301_),
    .Q(dbg_0.mem_data_12_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07037_ (
    .CLK(dco_clk),
    .D(_00302_),
    .Q(dbg_0.mem_data_13_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07038_ (
    .CLK(dco_clk),
    .D(_00303_),
    .Q(dbg_0.mem_data_14_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07039_ (
    .CLK(dco_clk),
    .D(_00304_),
    .Q(dbg_0.mem_data_15_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07040_ (
    .CLK(dco_clk),
    .D(_00314_),
    .Q(dbg_0.mem_start ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07041_ (
    .CLK(dco_clk),
    .D(_00295_),
    .Q(dbg_0.mem_ctl_1_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07042_ (
    .CLK(dco_clk),
    .D(_00296_),
    .Q(dbg_0.mem_ctl_2_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07043_ (
    .CLK(dco_clk),
    .D(_00297_),
    .Q(dbg_0.dbg_i2c_0.mem_bw ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07044_ (
    .CLK(dco_clk),
    .D(_00257_),
    .Q(dbg_0.cpu_stat_2_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07045_ (
    .CLK(dco_clk),
    .D(_00258_),
    .Q(dbg_0.cpu_stat_3_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07046_ (
    .CLK(dco_clk),
    .D(_00253_),
    .Q(dbg_0.cpu_ctl_3_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07047_ (
    .CLK(dco_clk),
    .D(_00254_),
    .Q(dbg_0.cpu_ctl_4_ ),
    .R(1'h1),
    .S(_00320_)
  );
  DFFSR _07048_ (
    .CLK(dco_clk),
    .D(_00255_),
    .Q(dbg_0.cpu_ctl_5_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07049_ (
    .CLK(dco_clk),
    .D(_00256_),
    .Q(clock_module_0.dbg_cpu_reset ),
    .R(_00320_),
    .S(1'h1)
  );
  INVX1 _07050_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_4_ ),
    .Y(_00821_)
  );
  INVX1 _07051_ (
    .A(dbg_0.dbg_i2c_0.sda_in_dly ),
    .Y(_00822_)
  );
  INVX1 _07052_ (
    .A(dbg_0.dbg_i2c_0.sda_in_sync_n ),
    .Y(dbg_0.dbg_i2c_0.sda_in_sync )
  );
  INVX1 _07053_ (
    .A(dbg_0.dbg_i2c_0.scl_sync_n ),
    .Y(dbg_0.dbg_i2c_0.scl_sync )
  );
  INVX1 _07054_ (
    .A(dbg_0.dbg_i2c_0.i2c_active_seq ),
    .Y(_00823_)
  );
  INVX1 _07055_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .Y(_00824_)
  );
  INVX1 _07056_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .Y(_00825_)
  );
  INVX1 _07057_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .Y(_00826_)
  );
  INVX1 _07058_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_4_ ),
    .Y(_00827_)
  );
  INVX1 _07059_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .Y(_00828_)
  );
  INVX1 _07060_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00829_)
  );
  INVX1 _07061_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .Y(_00830_)
  );
  INVX1 _07062_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .Y(_00831_)
  );
  INVX1 _07063_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_3_ ),
    .Y(_00832_)
  );
  INVX1 _07064_ (
    .A(dbg_0.dbg_din_8_ ),
    .Y(_00833_)
  );
  INVX1 _07065_ (
    .A(dbg_0.dbg_din_9_ ),
    .Y(_00834_)
  );
  INVX1 _07066_ (
    .A(dbg_0.dbg_din_10_ ),
    .Y(_00835_)
  );
  INVX1 _07067_ (
    .A(dbg_0.dbg_din_11_ ),
    .Y(_00836_)
  );
  INVX1 _07068_ (
    .A(dbg_0.dbg_din_12_ ),
    .Y(_00837_)
  );
  INVX1 _07069_ (
    .A(dbg_0.dbg_din_13_ ),
    .Y(_00838_)
  );
  INVX1 _07070_ (
    .A(dbg_0.dbg_din_14_ ),
    .Y(_00839_)
  );
  INVX1 _07071_ (
    .A(dbg_0.dbg_din_15_ ),
    .Y(_00840_)
  );
  INVX1 _07072_ (
    .A(dbg_0.dbg_dout_0_ ),
    .Y(_00841_)
  );
  INVX1 _07073_ (
    .A(dbg_0.dbg_dout_1_ ),
    .Y(_00842_)
  );
  INVX1 _07074_ (
    .A(dbg_0.dbg_dout_2_ ),
    .Y(_00843_)
  );
  INVX1 _07075_ (
    .A(dbg_0.dbg_dout_3_ ),
    .Y(_00844_)
  );
  INVX1 _07076_ (
    .A(dbg_0.dbg_dout_4_ ),
    .Y(_00845_)
  );
  INVX1 _07077_ (
    .A(dbg_0.dbg_dout_5_ ),
    .Y(_00846_)
  );
  INVX1 _07078_ (
    .A(dbg_0.dbg_dout_6_ ),
    .Y(_00847_)
  );
  INVX1 _07079_ (
    .A(dbg_0.dbg_dout_7_ ),
    .Y(_00848_)
  );
  INVX1 _07080_ (
    .A(dbg_i2c_scl),
    .Y(dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_in )
  );
  INVX1 _07081_ (
    .A(dbg_i2c_sda_in),
    .Y(dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_in )
  );
  INVX1 _07082_ (
    .A(clock_module_0.dbg_rst ),
    .Y(_00820_)
  );
  OR2X1 _07083_ (
    .A(dbg_0.dbg_i2c_0.sda_in_buf_1_ ),
    .B(dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .Y(_00849_)
  );
  AND2X1 _07084_ (
    .A(dbg_0.dbg_i2c_0.sda_in_buf_1_ ),
    .B(dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .Y(_00850_)
  );
  OAI21X1 _07085_ (
    .A(dbg_0.dbg_i2c_0.sda_in_sync ),
    .B(_00850_),
    .C(_00849_),
    .Y(_00851_)
  );
  INVX1 _07086_ (
    .A(_00851_),
    .Y(dbg_0.dbg_i2c_0.sda_in )
  );
  OR2X1 _07087_ (
    .A(dbg_0.dbg_i2c_0.scl_buf_1_ ),
    .B(dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .Y(_00852_)
  );
  AND2X1 _07088_ (
    .A(dbg_0.dbg_i2c_0.scl_buf_1_ ),
    .B(dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .Y(_00853_)
  );
  OAI21X1 _07089_ (
    .A(dbg_0.dbg_i2c_0.scl_sync ),
    .B(_00853_),
    .C(_00852_),
    .Y(_00854_)
  );
  INVX1 _07090_ (
    .A(_00854_),
    .Y(dbg_0.dbg_i2c_0.scl )
  );
  XNOR2X1 _07091_ (
    .A(dbg_i2c_addr_4_),
    .B(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .Y(_00855_)
  );
  XNOR2X1 _07092_ (
    .A(dbg_i2c_addr_2_),
    .B(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .Y(_00856_)
  );
  XNOR2X1 _07093_ (
    .A(dbg_i2c_addr_1_),
    .B(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .Y(_00857_)
  );
  NAND3X1 _07094_ (
    .A(_00855_),
    .B(_00856_),
    .C(_00857_),
    .Y(_00858_)
  );
  XNOR2X1 _07095_ (
    .A(dbg_i2c_addr_6_),
    .B(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .Y(_00859_)
  );
  XNOR2X1 _07096_ (
    .A(dbg_i2c_addr_0_),
    .B(dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .Y(_00860_)
  );
  XOR2X1 _07097_ (
    .A(dbg_i2c_addr_5_),
    .B(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .Y(_00861_)
  );
  XOR2X1 _07098_ (
    .A(dbg_i2c_addr_3_),
    .B(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .Y(_00862_)
  );
  NOR2X1 _07099_ (
    .A(_00861_),
    .B(_00862_),
    .Y(_00863_)
  );
  NAND3X1 _07100_ (
    .A(_00859_),
    .B(_00860_),
    .C(_00863_),
    .Y(_00864_)
  );
  NOR2X1 _07101_ (
    .A(_00858_),
    .B(_00864_),
    .Y(_00865_)
  );
  INVX1 _07102_ (
    .A(_00865_),
    .Y(_00866_)
  );
  AND2X1 _07103_ (
    .A(dbg_0.dbg_i2c_0.scl_dly ),
    .B(_00854_),
    .Y(_00867_)
  );
  NAND2X1 _07104_ (
    .A(dbg_0.dbg_i2c_0.scl_dly ),
    .B(_00854_),
    .Y(_00868_)
  );
  NAND2X1 _07105_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .B(_00867_),
    .Y(_00869_)
  );
  OAI21X1 _07106_ (
    .A(_00866_),
    .B(_00869_),
    .C(dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .Y(_00870_)
  );
  NOR3X1 _07107_ (
    .A(_00822_),
    .B(dbg_0.dbg_i2c_0.sda_in ),
    .C(_00854_),
    .Y(_00871_)
  );
  NAND3X1 _07108_ (
    .A(dbg_0.dbg_i2c_0.sda_in_dly ),
    .B(_00851_),
    .C(dbg_0.dbg_i2c_0.scl ),
    .Y(_00872_)
  );
  NOR3X1 _07109_ (
    .A(dbg_0.dbg_i2c_0.sda_in_dly ),
    .B(_00851_),
    .C(_00854_),
    .Y(_00873_)
  );
  NAND3X1 _07110_ (
    .A(_00822_),
    .B(dbg_0.dbg_i2c_0.sda_in ),
    .C(dbg_0.dbg_i2c_0.scl ),
    .Y(_00874_)
  );
  NOR2X1 _07111_ (
    .A(_00823_),
    .B(_00873_),
    .Y(_00875_)
  );
  NOR3X1 _07112_ (
    .A(_00823_),
    .B(_00871_),
    .C(_00873_),
    .Y(_00876_)
  );
  NAND3X1 _07113_ (
    .A(dbg_0.dbg_i2c_0.i2c_active_seq ),
    .B(_00872_),
    .C(_00874_),
    .Y(_00877_)
  );
  NAND3X1 _07114_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_4_ ),
    .B(dbg_0.dbg_i2c_0.sda_in ),
    .C(_00867_),
    .Y(_00878_)
  );
  NOR2X1 _07115_ (
    .A(_00825_),
    .B(_00869_),
    .Y(_00879_)
  );
  OR2X1 _07116_ (
    .A(_00825_),
    .B(_00869_),
    .Y(_00880_)
  );
  NAND3X1 _07117_ (
    .A(_00870_),
    .B(_00876_),
    .C(_00878_),
    .Y(_00814_)
  );
  NOR2X1 _07118_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .B(dbg_0.dbg_i2c_0.i2c_state_5_ ),
    .Y(_00881_)
  );
  NAND2X1 _07119_ (
    .A(_00825_),
    .B(_00881_),
    .Y(_00882_)
  );
  NOR2X1 _07120_ (
    .A(_00824_),
    .B(_00869_),
    .Y(_00883_)
  );
  OR2X1 _07121_ (
    .A(_00824_),
    .B(_00869_),
    .Y(_00884_)
  );
  NOR2X1 _07122_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .B(_00884_),
    .Y(_00885_)
  );
  NOR2X1 _07123_ (
    .A(_00831_),
    .B(dbg_0.dbg_i2c_0.mem_burst_wr ),
    .Y(_00886_)
  );
  OAI21X1 _07124_ (
    .A(dbg_0.dbg_i2c_0.mem_burst_rd ),
    .B(_00885_),
    .C(_00886_),
    .Y(_00887_)
  );
  AND2X1 _07125_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_i2c_0.mem_bw ),
    .Y(_00888_)
  );
  OR2X1 _07126_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .Y(_00889_)
  );
  NOR2X1 _07127_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00889_),
    .Y(_00890_)
  );
  OR2X1 _07128_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00889_),
    .Y(_00891_)
  );
  AND2X1 _07129_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .B(_00826_),
    .Y(_00892_)
  );
  NOR2X1 _07130_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .Y(_00893_)
  );
  NOR2X1 _07131_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .Y(_00894_)
  );
  AND2X1 _07132_ (
    .A(_00893_),
    .B(_00894_),
    .Y(_00895_)
  );
  NAND3X1 _07133_ (
    .A(_00890_),
    .B(_00892_),
    .C(_00895_),
    .Y(_00896_)
  );
  NOR2X1 _07134_ (
    .A(_00868_),
    .B(_00896_),
    .Y(_00897_)
  );
  OAI21X1 _07135_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_4_ ),
    .B(dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .C(_00897_),
    .Y(_00898_)
  );
  OR2X1 _07136_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .Y(_00899_)
  );
  NOR2X1 _07137_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .Y(_00900_)
  );
  NAND3X1 _07138_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .B(_00826_),
    .C(_00900_),
    .Y(_00901_)
  );
  NOR3X1 _07139_ (
    .A(_00891_),
    .B(_00899_),
    .C(_00901_),
    .Y(_00902_)
  );
  OAI21X1 _07140_ (
    .A(_00888_),
    .B(_00898_),
    .C(dbg_0.dbg_i2c_0.dbg_state_4_ ),
    .Y(_00903_)
  );
  NOR2X1 _07141_ (
    .A(_00830_),
    .B(_00898_),
    .Y(_00904_)
  );
  NAND2X1 _07142_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(_00904_),
    .Y(_00905_)
  );
  NAND3X1 _07143_ (
    .A(_00887_),
    .B(_00903_),
    .C(_00905_),
    .Y(_00813_)
  );
  NAND2X1 _07144_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(dbg_0.dbg_i2c_0.i2c_state_3_ ),
    .Y(_00906_)
  );
  NAND2X1 _07145_ (
    .A(_00821_),
    .B(_00906_),
    .Y(_00907_)
  );
  OAI21X1 _07146_ (
    .A(_00821_),
    .B(dbg_0.dbg_i2c_0.sda_in ),
    .C(_00906_),
    .Y(_00908_)
  );
  NAND2X1 _07147_ (
    .A(_00867_),
    .B(_00908_),
    .Y(_00909_)
  );
  OAI21X1 _07148_ (
    .A(_00868_),
    .B(_00896_),
    .C(dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .Y(_00910_)
  );
  AOI21X1 _07149_ (
    .A(_00909_),
    .B(_00910_),
    .C(_00877_),
    .Y(_00815_)
  );
  AND2X1 _07150_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00898_),
    .Y(_00911_)
  );
  AOI21X1 _07151_ (
    .A(_00829_),
    .B(dbg_0.dbg_i2c_0.dbg_bw ),
    .C(_00888_),
    .Y(_00912_)
  );
  NOR2X1 _07152_ (
    .A(_00827_),
    .B(_00898_),
    .Y(_00913_)
  );
  AND2X1 _07153_ (
    .A(_00912_),
    .B(_00913_),
    .Y(_00914_)
  );
  OR2X1 _07154_ (
    .A(_00911_),
    .B(_00914_),
    .Y(_00810_)
  );
  NAND2X1 _07155_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_3_ ),
    .B(_00883_),
    .Y(_00915_)
  );
  OAI21X1 _07156_ (
    .A(_00827_),
    .B(_00898_),
    .C(_00915_),
    .Y(_00916_)
  );
  NAND3X1 _07157_ (
    .A(_00829_),
    .B(dbg_0.dbg_i2c_0.dbg_bw ),
    .C(_00916_),
    .Y(_00917_)
  );
  NOR2X1 _07158_ (
    .A(_00829_),
    .B(dbg_0.dbg_i2c_0.mem_burst_end ),
    .Y(_00918_)
  );
  NAND2X1 _07159_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_2_ ),
    .B(_00883_),
    .Y(_00919_)
  );
  NOR2X1 _07160_ (
    .A(dbg_0.dbg_i2c_0.mem_burst_rd ),
    .B(dbg_0.dbg_i2c_0.mem_burst_wr ),
    .Y(_00920_)
  );
  AND2X1 _07161_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .B(_00920_),
    .Y(_00921_)
  );
  NAND2X1 _07162_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_i2c_0.mem_burst_end ),
    .Y(_00922_)
  );
  NOR2X1 _07163_ (
    .A(_00832_),
    .B(_00922_),
    .Y(_00923_)
  );
  AOI21X1 _07164_ (
    .A(_00884_),
    .B(_00921_),
    .C(_00923_),
    .Y(_00924_)
  );
  OAI21X1 _07165_ (
    .A(_00918_),
    .B(_00919_),
    .C(_00924_),
    .Y(_00925_)
  );
  AOI21X1 _07166_ (
    .A(_00829_),
    .B(_00904_),
    .C(_00925_),
    .Y(_00926_)
  );
  NAND2X1 _07167_ (
    .A(_00917_),
    .B(_00926_),
    .Y(_00809_)
  );
  OAI21X1 _07168_ (
    .A(_00884_),
    .B(_00888_),
    .C(dbg_0.dbg_i2c_0.dbg_state_3_ ),
    .Y(_00927_)
  );
  OAI21X1 _07169_ (
    .A(_00829_),
    .B(_00919_),
    .C(_00927_),
    .Y(_00928_)
  );
  NOR2X1 _07170_ (
    .A(_00831_),
    .B(_00884_),
    .Y(_00929_)
  );
  NAND2X1 _07171_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .B(_00883_),
    .Y(_00930_)
  );
  NAND2X1 _07172_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .B(_00920_),
    .Y(_00931_)
  );
  AOI22X1 _07173_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .B(dbg_0.dbg_i2c_0.mem_burst_wr ),
    .C(_00922_),
    .D(_00928_),
    .Y(_00932_)
  );
  OAI21X1 _07174_ (
    .A(_00930_),
    .B(_00931_),
    .C(_00932_),
    .Y(_00812_)
  );
  OAI21X1 _07175_ (
    .A(_00824_),
    .B(_00869_),
    .C(dbg_0.dbg_i2c_0.dbg_state_2_ ),
    .Y(_00933_)
  );
  OAI21X1 _07176_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_i2c_0.dbg_bw ),
    .C(dbg_0.dbg_i2c_0.mem_burst_end ),
    .Y(_00934_)
  );
  NAND2X1 _07177_ (
    .A(_00912_),
    .B(_00934_),
    .Y(_00935_)
  );
  OAI21X1 _07178_ (
    .A(_00915_),
    .B(_00935_),
    .C(_00933_),
    .Y(_00811_)
  );
  NAND2X1 _07179_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_4_ ),
    .B(_00868_),
    .Y(_00936_)
  );
  NAND3X1 _07180_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .B(_00867_),
    .C(_00902_),
    .Y(_00937_)
  );
  NOR2X1 _07181_ (
    .A(_00867_),
    .B(_00877_),
    .Y(_00938_)
  );
  AOI21X1 _07182_ (
    .A(_00936_),
    .B(_00937_),
    .C(_00877_),
    .Y(_00818_)
  );
  NAND2X1 _07183_ (
    .A(_00876_),
    .B(_00883_),
    .Y(_00939_)
  );
  NAND2X1 _07184_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_5_ ),
    .B(_00938_),
    .Y(_00940_)
  );
  OAI21X1 _07185_ (
    .A(_00877_),
    .B(_00884_),
    .C(_00940_),
    .Y(_00819_)
  );
  NAND2X1 _07186_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_3_ ),
    .B(_00938_),
    .Y(_00941_)
  );
  NAND3X1 _07187_ (
    .A(_00865_),
    .B(_00876_),
    .C(_00879_),
    .Y(_00942_)
  );
  NAND2X1 _07188_ (
    .A(_00941_),
    .B(_00942_),
    .Y(_00817_)
  );
  NAND2X1 _07189_ (
    .A(_00828_),
    .B(dbg_0.dbg_i2c_0.i2c_state_3_ ),
    .Y(_00943_)
  );
  NAND2X1 _07190_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_5_ ),
    .B(_00867_),
    .Y(_00944_)
  );
  OAI21X1 _07191_ (
    .A(_00868_),
    .B(_00943_),
    .C(_00944_),
    .Y(_00945_)
  );
  AOI21X1 _07192_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .B(_00869_),
    .C(_00945_),
    .Y(_00946_)
  );
  NOR2X1 _07193_ (
    .A(_00877_),
    .B(_00946_),
    .Y(_00816_)
  );
  NOR2X1 _07194_ (
    .A(_00815_),
    .B(_00818_),
    .Y(_00947_)
  );
  OR2X1 _07195_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_5_ ),
    .B(dbg_0.dbg_i2c_0.i2c_state_3_ ),
    .Y(_00948_)
  );
  OAI21X1 _07196_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_4_ ),
    .B(_00948_),
    .C(_00938_),
    .Y(_00949_)
  );
  NAND3X1 _07197_ (
    .A(_00939_),
    .B(_00942_),
    .C(_00949_),
    .Y(_00950_)
  );
  AND2X1 _07198_ (
    .A(_00947_),
    .B(_00950_),
    .Y(_00951_)
  );
  OAI21X1 _07199_ (
    .A(_00868_),
    .B(_00943_),
    .C(_00881_),
    .Y(_00952_)
  );
  NAND2X1 _07200_ (
    .A(_00867_),
    .B(_00896_),
    .Y(_00953_)
  );
  AOI21X1 _07201_ (
    .A(_00876_),
    .B(_00952_),
    .C(_00953_),
    .Y(_00954_)
  );
  OAI21X1 _07202_ (
    .A(_00815_),
    .B(_00818_),
    .C(_00954_),
    .Y(_00955_)
  );
  NAND2X1 _07203_ (
    .A(_00050_),
    .B(_00868_),
    .Y(_00956_)
  );
  OAI21X1 _07204_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .B(_00955_),
    .C(_00867_),
    .Y(_00957_)
  );
  OAI21X1 _07205_ (
    .A(_00951_),
    .B(_00957_),
    .C(_00956_),
    .Y(_00805_)
  );
  MUX2X1 _07206_ (
    .A(dbg_0.dbg_din_0_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .S(_00915_),
    .Y(_00958_)
  );
  INVX1 _07207_ (
    .A(_00958_),
    .Y(_00797_)
  );
  MUX2X1 _07208_ (
    .A(dbg_0.dbg_din_1_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .S(_00915_),
    .Y(_00959_)
  );
  INVX1 _07209_ (
    .A(_00959_),
    .Y(_00798_)
  );
  MUX2X1 _07210_ (
    .A(dbg_0.dbg_din_2_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .S(_00915_),
    .Y(_00960_)
  );
  INVX1 _07211_ (
    .A(_00960_),
    .Y(_00799_)
  );
  MUX2X1 _07212_ (
    .A(dbg_0.dbg_din_3_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .S(_00915_),
    .Y(_00961_)
  );
  INVX1 _07213_ (
    .A(_00961_),
    .Y(_00800_)
  );
  MUX2X1 _07214_ (
    .A(dbg_0.dbg_din_4_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .S(_00915_),
    .Y(_00962_)
  );
  INVX1 _07215_ (
    .A(_00962_),
    .Y(_00801_)
  );
  MUX2X1 _07216_ (
    .A(dbg_0.dbg_din_5_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .S(_00915_),
    .Y(_00963_)
  );
  INVX1 _07217_ (
    .A(_00963_),
    .Y(_00802_)
  );
  MUX2X1 _07218_ (
    .A(dbg_0.dbg_din_6_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .S(_00915_),
    .Y(_00964_)
  );
  INVX1 _07219_ (
    .A(_00964_),
    .Y(_00803_)
  );
  MUX2X1 _07220_ (
    .A(dbg_0.dbg_din_7_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .S(_00915_),
    .Y(_00965_)
  );
  INVX1 _07221_ (
    .A(_00965_),
    .Y(_00804_)
  );
  NAND3X1 _07222_ (
    .A(_00829_),
    .B(dbg_0.dbg_addr_0_ ),
    .C(_00930_),
    .Y(_00966_)
  );
  OAI21X1 _07223_ (
    .A(_00828_),
    .B(_00930_),
    .C(_00966_),
    .Y(_00782_)
  );
  OAI21X1 _07224_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_addr_1_ ),
    .C(_00930_),
    .Y(_00967_)
  );
  OAI21X1 _07225_ (
    .A(_00826_),
    .B(_00930_),
    .C(_00967_),
    .Y(_00783_)
  );
  NOR2X1 _07226_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_addr_2_ ),
    .Y(_00968_)
  );
  NAND2X1 _07227_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B(_00929_),
    .Y(_00969_)
  );
  OAI21X1 _07228_ (
    .A(_00929_),
    .B(_00968_),
    .C(_00969_),
    .Y(_00784_)
  );
  NAND2X1 _07229_ (
    .A(_00829_),
    .B(dbg_0.dbg_addr_3_ ),
    .Y(_00970_)
  );
  NAND2X1 _07230_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .B(_00929_),
    .Y(_00971_)
  );
  OAI21X1 _07231_ (
    .A(_00929_),
    .B(_00970_),
    .C(_00971_),
    .Y(_00785_)
  );
  NAND2X1 _07232_ (
    .A(_00829_),
    .B(dbg_0.dbg_addr_4_ ),
    .Y(_00972_)
  );
  NAND2X1 _07233_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B(_00929_),
    .Y(_00973_)
  );
  OAI21X1 _07234_ (
    .A(_00929_),
    .B(_00972_),
    .C(_00973_),
    .Y(_00786_)
  );
  NAND2X1 _07235_ (
    .A(_00829_),
    .B(dbg_0.dbg_addr_5_ ),
    .Y(_00974_)
  );
  NAND2X1 _07236_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .B(_00929_),
    .Y(_00975_)
  );
  OAI21X1 _07237_ (
    .A(_00929_),
    .B(_00974_),
    .C(_00975_),
    .Y(_00787_)
  );
  NAND2X1 _07238_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(_00929_),
    .Y(_00976_)
  );
  OAI21X1 _07239_ (
    .A(_00912_),
    .B(_00929_),
    .C(_00976_),
    .Y(_00788_)
  );
  OAI21X1 _07240_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00919_),
    .C(_00915_),
    .Y(_00977_)
  );
  AOI21X1 _07241_ (
    .A(_00833_),
    .B(_00919_),
    .C(_00977_),
    .Y(_00789_)
  );
  OAI21X1 _07242_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .B(_00919_),
    .C(_00915_),
    .Y(_00978_)
  );
  AOI21X1 _07243_ (
    .A(_00834_),
    .B(_00919_),
    .C(_00978_),
    .Y(_00790_)
  );
  OAI21X1 _07244_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B(_00919_),
    .C(_00915_),
    .Y(_00979_)
  );
  AOI21X1 _07245_ (
    .A(_00835_),
    .B(_00919_),
    .C(_00979_),
    .Y(_00791_)
  );
  OAI21X1 _07246_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .B(_00919_),
    .C(_00915_),
    .Y(_00980_)
  );
  AOI21X1 _07247_ (
    .A(_00836_),
    .B(_00919_),
    .C(_00980_),
    .Y(_00792_)
  );
  OAI21X1 _07248_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B(_00919_),
    .C(_00915_),
    .Y(_00981_)
  );
  AOI21X1 _07249_ (
    .A(_00837_),
    .B(_00919_),
    .C(_00981_),
    .Y(_00793_)
  );
  OAI21X1 _07250_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .B(_00919_),
    .C(_00915_),
    .Y(_00982_)
  );
  AOI21X1 _07251_ (
    .A(_00838_),
    .B(_00919_),
    .C(_00982_),
    .Y(_00794_)
  );
  OAI21X1 _07252_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(_00919_),
    .C(_00915_),
    .Y(_00983_)
  );
  AOI21X1 _07253_ (
    .A(_00839_),
    .B(_00919_),
    .C(_00983_),
    .Y(_00795_)
  );
  OAI21X1 _07254_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .B(_00919_),
    .C(_00915_),
    .Y(_00984_)
  );
  AOI21X1 _07255_ (
    .A(_00840_),
    .B(_00919_),
    .C(_00984_),
    .Y(_00796_)
  );
  NOR2X1 _07256_ (
    .A(dbg_0.dbg_i2c_0.scl_dly ),
    .B(_00854_),
    .Y(dbg_0.dbg_i2c_0.scl_re )
  );
  NAND2X1 _07257_ (
    .A(dbg_0.dbg_i2c_0.scl_re_dly_1_ ),
    .B(_00882_),
    .Y(_00985_)
  );
  NAND2X1 _07258_ (
    .A(_00955_),
    .B(_00985_),
    .Y(_00986_)
  );
  NOR2X1 _07259_ (
    .A(_00877_),
    .B(_00945_),
    .Y(_00987_)
  );
  NAND2X1 _07260_ (
    .A(_00907_),
    .B(dbg_0.dbg_i2c_0.scl_re ),
    .Y(_00988_)
  );
  OAI21X1 _07261_ (
    .A(_00851_),
    .B(_00985_),
    .C(_00987_),
    .Y(_00989_)
  );
  AOI21X1 _07262_ (
    .A(_00907_),
    .B(dbg_0.dbg_i2c_0.scl_re ),
    .C(_00989_),
    .Y(_00990_)
  );
  OAI21X1 _07263_ (
    .A(_00828_),
    .B(_00986_),
    .C(_00990_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_0_ )
  );
  MUX2X1 _07264_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .S(_00986_),
    .Y(_00991_)
  );
  NAND2X1 _07265_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_8_ ),
    .Y(_00992_)
  );
  OAI21X1 _07266_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00841_),
    .C(_00992_),
    .Y(_00993_)
  );
  OAI21X1 _07267_ (
    .A(_00988_),
    .B(_00993_),
    .C(_00987_),
    .Y(_00994_)
  );
  AOI21X1 _07268_ (
    .A(_00988_),
    .B(_00991_),
    .C(_00994_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_1_ )
  );
  MUX2X1 _07269_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .S(_00986_),
    .Y(_00995_)
  );
  NAND2X1 _07270_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_9_ ),
    .Y(_00996_)
  );
  OAI21X1 _07271_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00842_),
    .C(_00996_),
    .Y(_00997_)
  );
  OAI21X1 _07272_ (
    .A(_00988_),
    .B(_00997_),
    .C(_00987_),
    .Y(_00998_)
  );
  AOI21X1 _07273_ (
    .A(_00988_),
    .B(_00995_),
    .C(_00998_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_2_ )
  );
  MUX2X1 _07274_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .S(_00986_),
    .Y(_00999_)
  );
  NAND2X1 _07275_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_10_ ),
    .Y(_01000_)
  );
  OAI21X1 _07276_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00843_),
    .C(_01000_),
    .Y(_01001_)
  );
  OAI21X1 _07277_ (
    .A(_00988_),
    .B(_01001_),
    .C(_00987_),
    .Y(_01002_)
  );
  AOI21X1 _07278_ (
    .A(_00988_),
    .B(_00999_),
    .C(_01002_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_3_ )
  );
  MUX2X1 _07279_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .S(_00986_),
    .Y(_01003_)
  );
  NAND2X1 _07280_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_11_ ),
    .Y(_01004_)
  );
  OAI21X1 _07281_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00844_),
    .C(_01004_),
    .Y(_01005_)
  );
  OAI21X1 _07282_ (
    .A(_00988_),
    .B(_01005_),
    .C(_00987_),
    .Y(_01006_)
  );
  AOI21X1 _07283_ (
    .A(_00988_),
    .B(_01003_),
    .C(_01006_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_4_ )
  );
  MUX2X1 _07284_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .S(_00986_),
    .Y(_01007_)
  );
  NAND2X1 _07285_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_12_ ),
    .Y(_01008_)
  );
  OAI21X1 _07286_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00845_),
    .C(_01008_),
    .Y(_01009_)
  );
  OAI21X1 _07287_ (
    .A(_00988_),
    .B(_01009_),
    .C(_00987_),
    .Y(_01010_)
  );
  AOI21X1 _07288_ (
    .A(_00988_),
    .B(_01007_),
    .C(_01010_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_5_ )
  );
  MUX2X1 _07289_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .S(_00986_),
    .Y(_01011_)
  );
  NAND2X1 _07290_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_13_ ),
    .Y(_01012_)
  );
  OAI21X1 _07291_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00846_),
    .C(_01012_),
    .Y(_01013_)
  );
  OAI21X1 _07292_ (
    .A(_00988_),
    .B(_01013_),
    .C(_00987_),
    .Y(_01014_)
  );
  AOI21X1 _07293_ (
    .A(_00988_),
    .B(_01011_),
    .C(_01014_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_6_ )
  );
  MUX2X1 _07294_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .S(_00986_),
    .Y(_01015_)
  );
  NAND2X1 _07295_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_14_ ),
    .Y(_01016_)
  );
  OAI21X1 _07296_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00847_),
    .C(_01016_),
    .Y(_01017_)
  );
  OAI21X1 _07297_ (
    .A(_00988_),
    .B(_01017_),
    .C(_00987_),
    .Y(_01018_)
  );
  AOI21X1 _07298_ (
    .A(_00988_),
    .B(_01015_),
    .C(_01018_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_7_ )
  );
  MUX2X1 _07299_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .S(_00986_),
    .Y(_01019_)
  );
  NAND2X1 _07300_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_15_ ),
    .Y(_01020_)
  );
  OAI21X1 _07301_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00848_),
    .C(_01020_),
    .Y(_01021_)
  );
  OAI21X1 _07302_ (
    .A(_00988_),
    .B(_01021_),
    .C(_00987_),
    .Y(_01022_)
  );
  AOI21X1 _07303_ (
    .A(_00988_),
    .B(_01019_),
    .C(_01022_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_8_ )
  );
  MUX2X1 _07304_ (
    .A(_00919_),
    .B(_00915_),
    .S(_00912_),
    .Y(_00807_)
  );
  NOR2X1 _07305_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .B(dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_01023_)
  );
  AOI22X1 _07306_ (
    .A(_00888_),
    .B(_00913_),
    .C(_00929_),
    .D(_01023_),
    .Y(_01024_)
  );
  OAI21X1 _07307_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00905_),
    .C(_01024_),
    .Y(_00806_)
  );
  OAI21X1 _07308_ (
    .A(_00865_),
    .B(_00880_),
    .C(_00875_),
    .Y(_01025_)
  );
  NAND2X1 _07309_ (
    .A(_00872_),
    .B(_01025_),
    .Y(_00808_)
  );
  DFFSR _07310_ (
    .CLK(dco_clk),
    .D(_00814_),
    .Q(dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .R(1'h1),
    .S(_00820_)
  );
  DFFSR _07311_ (
    .CLK(dco_clk),
    .D(_00815_),
    .Q(dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07312_ (
    .CLK(dco_clk),
    .D(_00816_),
    .Q(dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07313_ (
    .CLK(dco_clk),
    .D(_00817_),
    .Q(dbg_0.dbg_i2c_0.i2c_state_3_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07314_ (
    .CLK(dco_clk),
    .D(_00818_),
    .Q(dbg_0.dbg_i2c_0.i2c_state_4_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07315_ (
    .CLK(dco_clk),
    .D(_00819_),
    .Q(dbg_0.dbg_i2c_0.i2c_state_5_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07316_ (
    .CLK(dco_clk),
    .D(_00809_),
    .Q(dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .R(1'h1),
    .S(_00820_)
  );
  DFFSR _07317_ (
    .CLK(dco_clk),
    .D(_00810_),
    .Q(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07318_ (
    .CLK(dco_clk),
    .D(_00811_),
    .Q(dbg_0.dbg_i2c_0.dbg_state_2_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07319_ (
    .CLK(dco_clk),
    .D(_00812_),
    .Q(dbg_0.dbg_i2c_0.dbg_state_3_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07320_ (
    .CLK(dco_clk),
    .D(_00813_),
    .Q(dbg_0.dbg_i2c_0.dbg_state_4_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07321_ (
    .CLK(dco_clk),
    .D(_00806_),
    .Q(dbg_0.dbg_i2c_0.dbg_rd ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07322_ (
    .CLK(dco_clk),
    .D(_00807_),
    .Q(dbg_0.dbg_i2c_0.dbg_wr ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07323_ (
    .CLK(dco_clk),
    .D(_00789_),
    .Q(dbg_0.dbg_din_8_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07324_ (
    .CLK(dco_clk),
    .D(_00790_),
    .Q(dbg_0.dbg_din_9_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07325_ (
    .CLK(dco_clk),
    .D(_00791_),
    .Q(dbg_0.dbg_din_10_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07326_ (
    .CLK(dco_clk),
    .D(_00792_),
    .Q(dbg_0.dbg_din_11_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07327_ (
    .CLK(dco_clk),
    .D(_00793_),
    .Q(dbg_0.dbg_din_12_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07328_ (
    .CLK(dco_clk),
    .D(_00794_),
    .Q(dbg_0.dbg_din_13_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07329_ (
    .CLK(dco_clk),
    .D(_00795_),
    .Q(dbg_0.dbg_din_14_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07330_ (
    .CLK(dco_clk),
    .D(_00796_),
    .Q(dbg_0.dbg_din_15_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07331_ (
    .CLK(dco_clk),
    .D(_00797_),
    .Q(dbg_0.dbg_din_0_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07332_ (
    .CLK(dco_clk),
    .D(_00798_),
    .Q(dbg_0.dbg_din_1_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07333_ (
    .CLK(dco_clk),
    .D(_00799_),
    .Q(dbg_0.dbg_din_2_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07334_ (
    .CLK(dco_clk),
    .D(_00800_),
    .Q(dbg_0.dbg_din_3_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07335_ (
    .CLK(dco_clk),
    .D(_00801_),
    .Q(dbg_0.dbg_din_4_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07336_ (
    .CLK(dco_clk),
    .D(_00802_),
    .Q(dbg_0.dbg_din_5_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07337_ (
    .CLK(dco_clk),
    .D(_00803_),
    .Q(dbg_0.dbg_din_6_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07338_ (
    .CLK(dco_clk),
    .D(_00804_),
    .Q(dbg_0.dbg_din_7_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07339_ (
    .CLK(dco_clk),
    .D(_00782_),
    .Q(dbg_0.dbg_addr_0_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07340_ (
    .CLK(dco_clk),
    .D(_00783_),
    .Q(dbg_0.dbg_addr_1_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07341_ (
    .CLK(dco_clk),
    .D(_00784_),
    .Q(dbg_0.dbg_addr_2_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07342_ (
    .CLK(dco_clk),
    .D(_00785_),
    .Q(dbg_0.dbg_addr_3_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07343_ (
    .CLK(dco_clk),
    .D(_00786_),
    .Q(dbg_0.dbg_addr_4_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07344_ (
    .CLK(dco_clk),
    .D(_00787_),
    .Q(dbg_0.dbg_addr_5_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07345_ (
    .CLK(dco_clk),
    .D(_00788_),
    .Q(dbg_0.dbg_i2c_0.dbg_bw ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07346_ (
    .CLK(dco_clk),
    .D(_00805_),
    .Q(_00050_),
    .R(1'h1),
    .S(_00820_)
  );
  DFFSR _07347_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_0_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .R(1'h1),
    .S(_00820_)
  );
  DFFSR _07348_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_1_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07349_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_2_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07350_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_3_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07351_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_4_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07352_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_5_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07353_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_6_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07354_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_7_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07355_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_8_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07356_ (
    .CLK(dco_clk),
    .D(_00808_),
    .Q(dbg_0.dbg_i2c_0.i2c_active_seq ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07357_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.scl_re ),
    .Q(dbg_0.dbg_i2c_0.scl_re_dly_0_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07358_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.scl_re_dly_0_ ),
    .Q(dbg_0.dbg_i2c_0.scl_re_dly_1_ ),
    .R(_00820_),
    .S(1'h1)
  );
  DFFSR _07359_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.scl ),
    .Q(dbg_0.dbg_i2c_0.scl_dly ),
    .R(1'h1),
    .S(_00820_)
  );
  DFFSR _07360_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.sda_in ),
    .Q(dbg_0.dbg_i2c_0.sda_in_dly ),
    .R(1'h1),
    .S(_00820_)
  );
  DFFSR _07361_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.sda_in_sync ),
    .Q(dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .R(1'h1),
    .S(_00820_)
  );
  DFFSR _07362_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .Q(dbg_0.dbg_i2c_0.sda_in_buf_1_ ),
    .R(1'h1),
    .S(_00820_)
  );
  DFFSR _07363_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.scl_sync ),
    .Q(dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .R(1'h1),
    .S(_00820_)
  );
  DFFSR _07364_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .Q(dbg_0.dbg_i2c_0.scl_buf_1_ ),
    .R(1'h1),
    .S(_00820_)
  );
  INVX1 _07365_ (
    .A(clock_module_0.dbg_rst ),
    .Y(_01026_)
  );
  DFFSR _07366_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_in ),
    .Q(dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_sync_0_ ),
    .R(_01026_),
    .S(1'h1)
  );
  DFFSR _07367_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_sync_0_ ),
    .Q(dbg_0.dbg_i2c_0.scl_sync_n ),
    .R(_01026_),
    .S(1'h1)
  );
  INVX1 _07368_ (
    .A(clock_module_0.dbg_rst ),
    .Y(_01027_)
  );
  DFFSR _07369_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_in ),
    .Q(dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_sync_0_ ),
    .R(_01027_),
    .S(1'h1)
  );
  DFFSR _07370_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_sync_0_ ),
    .Q(dbg_0.dbg_i2c_0.sda_in_sync_n ),
    .R(_01027_),
    .S(1'h1)
  );
  INVX1 _07371_ (
    .A(e_state_0_),
    .Y(_01064_)
  );
  INVX1 _07372_ (
    .A(e_state_2_),
    .Y(_01065_)
  );
  INVX1 _07373_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .Y(_01066_)
  );
  INVX1 _07374_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_alu ),
    .Y(_01067_)
  );
  INVX1 _07375_ (
    .A(execution_unit_0.mab_lsb ),
    .Y(_01068_)
  );
  INVX1 _07376_ (
    .A(dbg_0.UNUSED_eu_mab_0_ ),
    .Y(_01069_)
  );
  INVX1 _07377_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .Y(_01070_)
  );
  INVX1 _07378_ (
    .A(execution_unit_0.mdb_out_nxt_8_ ),
    .Y(_01071_)
  );
  INVX1 _07379_ (
    .A(execution_unit_0.mdb_out_nxt_9_ ),
    .Y(_01072_)
  );
  INVX1 _07380_ (
    .A(execution_unit_0.mdb_out_nxt_10_ ),
    .Y(_01073_)
  );
  INVX1 _07381_ (
    .A(execution_unit_0.mdb_out_nxt_11_ ),
    .Y(_01074_)
  );
  INVX1 _07382_ (
    .A(execution_unit_0.mdb_out_nxt_12_ ),
    .Y(_01075_)
  );
  INVX1 _07383_ (
    .A(execution_unit_0.mdb_out_nxt_13_ ),
    .Y(_01076_)
  );
  INVX1 _07384_ (
    .A(execution_unit_0.mdb_out_nxt_14_ ),
    .Y(_01077_)
  );
  INVX1 _07385_ (
    .A(execution_unit_0.mdb_out_nxt_15_ ),
    .Y(_01078_)
  );
  INVX1 _07386_ (
    .A(dbg_0.dbg_reg_din_1_ ),
    .Y(_01079_)
  );
  INVX1 _07387_ (
    .A(dbg_0.dbg_reg_din_2_ ),
    .Y(_01080_)
  );
  INVX1 _07388_ (
    .A(dbg_0.dbg_reg_din_3_ ),
    .Y(_01081_)
  );
  INVX1 _07389_ (
    .A(dbg_0.dbg_reg_din_4_ ),
    .Y(_01082_)
  );
  INVX1 _07390_ (
    .A(dbg_0.dbg_reg_din_5_ ),
    .Y(_01083_)
  );
  INVX1 _07391_ (
    .A(dbg_0.dbg_reg_din_6_ ),
    .Y(_01084_)
  );
  INVX1 _07392_ (
    .A(dbg_0.dbg_reg_din_7_ ),
    .Y(_01085_)
  );
  INVX1 _07393_ (
    .A(execution_unit_0.mdb_in_buf_8_ ),
    .Y(_01086_)
  );
  INVX1 _07394_ (
    .A(dbg_0.dbg_reg_din_8_ ),
    .Y(_01087_)
  );
  INVX1 _07395_ (
    .A(execution_unit_0.mdb_in_buf_9_ ),
    .Y(_01088_)
  );
  INVX1 _07396_ (
    .A(dbg_0.dbg_reg_din_9_ ),
    .Y(_01089_)
  );
  INVX1 _07397_ (
    .A(execution_unit_0.mdb_in_buf_10_ ),
    .Y(_01090_)
  );
  INVX1 _07398_ (
    .A(dbg_0.dbg_reg_din_10_ ),
    .Y(_01091_)
  );
  INVX1 _07399_ (
    .A(execution_unit_0.mdb_in_buf_11_ ),
    .Y(_01092_)
  );
  INVX1 _07400_ (
    .A(dbg_0.dbg_reg_din_11_ ),
    .Y(_01093_)
  );
  INVX1 _07401_ (
    .A(execution_unit_0.mdb_in_buf_12_ ),
    .Y(_01094_)
  );
  INVX1 _07402_ (
    .A(dbg_0.dbg_reg_din_12_ ),
    .Y(_01095_)
  );
  INVX1 _07403_ (
    .A(execution_unit_0.mdb_in_buf_13_ ),
    .Y(_01096_)
  );
  INVX1 _07404_ (
    .A(dbg_0.dbg_reg_din_13_ ),
    .Y(_01097_)
  );
  INVX1 _07405_ (
    .A(execution_unit_0.mdb_in_buf_14_ ),
    .Y(_01098_)
  );
  INVX1 _07406_ (
    .A(dbg_0.dbg_reg_din_14_ ),
    .Y(_01099_)
  );
  INVX1 _07407_ (
    .A(execution_unit_0.mdb_in_buf_15_ ),
    .Y(_01100_)
  );
  INVX1 _07408_ (
    .A(dbg_0.dbg_reg_din_15_ ),
    .Y(_01101_)
  );
  INVX1 _07409_ (
    .A(cpu_halt_st),
    .Y(_01102_)
  );
  INVX1 _07410_ (
    .A(dbg_0.dbg_reg_wr ),
    .Y(_01103_)
  );
  INVX1 _07411_ (
    .A(_00162_),
    .Y(_01063_)
  );
  AND2X1 _07412_ (
    .A(_01065_),
    .B(e_state_3_),
    .Y(_01104_)
  );
  AND2X1 _07413_ (
    .A(e_state_0_),
    .B(e_state_1_),
    .Y(_01105_)
  );
  NAND3X1 _07414_ (
    .A(_01065_),
    .B(e_state_3_),
    .C(_01105_),
    .Y(_01106_)
  );
  INVX1 _07415_ (
    .A(_01106_),
    .Y(execution_unit_0.alu_0.exec_cycle )
  );
  NOR2X1 _07416_ (
    .A(_01065_),
    .B(e_state_3_),
    .Y(_01107_)
  );
  NAND2X1 _07417_ (
    .A(e_state_1_),
    .B(_01107_),
    .Y(_01108_)
  );
  AND2X1 _07418_ (
    .A(_01064_),
    .B(e_state_1_),
    .Y(_01109_)
  );
  NAND2X1 _07419_ (
    .A(_01107_),
    .B(_01109_),
    .Y(_01110_)
  );
  INVX1 _07420_ (
    .A(_01110_),
    .Y(_01045_)
  );
  NOR2X1 _07421_ (
    .A(e_state_2_),
    .B(e_state_3_),
    .Y(_01111_)
  );
  NAND2X1 _07422_ (
    .A(_01064_),
    .B(_01111_),
    .Y(_01112_)
  );
  NOR2X1 _07423_ (
    .A(e_state_1_),
    .B(_01112_),
    .Y(execution_unit_0.reg_sr_clr )
  );
  NAND2X1 _07424_ (
    .A(e_state_0_),
    .B(_01111_),
    .Y(_01113_)
  );
  NOR2X1 _07425_ (
    .A(execution_unit_0.inst_irq_rst ),
    .B(_01113_),
    .Y(_01114_)
  );
  NAND2X1 _07426_ (
    .A(_01105_),
    .B(_01107_),
    .Y(_01115_)
  );
  NAND2X1 _07427_ (
    .A(_01104_),
    .B(_01109_),
    .Y(_01116_)
  );
  NAND3X1 _07428_ (
    .A(_01066_),
    .B(_01104_),
    .C(_01109_),
    .Y(_01117_)
  );
  OAI21X1 _07429_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01116_),
    .C(_01115_),
    .Y(_01118_)
  );
  OAI21X1 _07430_ (
    .A(_01114_),
    .B(_01118_),
    .C(_01067_),
    .Y(_01119_)
  );
  NOR2X1 _07431_ (
    .A(_01064_),
    .B(e_state_1_),
    .Y(_01120_)
  );
  AND2X1 _07432_ (
    .A(_01104_),
    .B(_01120_),
    .Y(_01121_)
  );
  NAND2X1 _07433_ (
    .A(_01104_),
    .B(_01120_),
    .Y(_01122_)
  );
  NOR2X1 _07434_ (
    .A(execution_unit_0.inst_type_0_ ),
    .B(execution_unit_0.inst_mov ),
    .Y(_01123_)
  );
  NAND2X1 _07435_ (
    .A(_01121_),
    .B(_01123_),
    .Y(_01124_)
  );
  OAI21X1 _07436_ (
    .A(execution_unit_0.inst_as_5_ ),
    .B(_01110_),
    .C(_01124_),
    .Y(_01125_)
  );
  AOI21X1 _07437_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(execution_unit_0.alu_0.exec_cycle ),
    .C(_01125_),
    .Y(_01126_)
  );
  NAND2X1 _07438_ (
    .A(_01119_),
    .B(_01126_),
    .Y(dbg_0.UNUSED_eu_mb_en )
  );
  MUX2X1 _07439_ (
    .A(_01069_),
    .B(_01068_),
    .S(dbg_0.UNUSED_eu_mb_en ),
    .Y(_01028_)
  );
  OAI21X1 _07440_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B(_01106_),
    .C(_01112_),
    .Y(_01127_)
  );
  MUX2X1 _07441_ (
    .A(execution_unit_0.alu_0.alu_out_0_ ),
    .B(eu_mdb_out_0_),
    .S(_01127_),
    .Y(_01128_)
  );
  NAND2X1 _07442_ (
    .A(UNUSED_fe_mab_0),
    .B(_01121_),
    .Y(_01129_)
  );
  OAI21X1 _07443_ (
    .A(_01121_),
    .B(_01128_),
    .C(_01129_),
    .Y(_01047_)
  );
  MUX2X1 _07444_ (
    .A(execution_unit_0.alu_0.alu_out_1_ ),
    .B(eu_mdb_out_1_),
    .S(_01127_),
    .Y(_01130_)
  );
  NAND2X1 _07445_ (
    .A(execution_unit_0.pc_nxt_1_ ),
    .B(_01121_),
    .Y(_01131_)
  );
  OAI21X1 _07446_ (
    .A(_01121_),
    .B(_01130_),
    .C(_01131_),
    .Y(_01054_)
  );
  MUX2X1 _07447_ (
    .A(execution_unit_0.alu_0.alu_out_2_ ),
    .B(eu_mdb_out_2_),
    .S(_01127_),
    .Y(_01132_)
  );
  NAND2X1 _07448_ (
    .A(execution_unit_0.pc_nxt_2_ ),
    .B(_01121_),
    .Y(_01133_)
  );
  OAI21X1 _07449_ (
    .A(_01121_),
    .B(_01132_),
    .C(_01133_),
    .Y(_01055_)
  );
  MUX2X1 _07450_ (
    .A(execution_unit_0.alu_0.alu_out_3_ ),
    .B(eu_mdb_out_3_),
    .S(_01127_),
    .Y(_01134_)
  );
  NAND2X1 _07451_ (
    .A(execution_unit_0.pc_nxt_3_ ),
    .B(_01121_),
    .Y(_01135_)
  );
  OAI21X1 _07452_ (
    .A(_01121_),
    .B(_01134_),
    .C(_01135_),
    .Y(_01056_)
  );
  MUX2X1 _07453_ (
    .A(execution_unit_0.alu_0.alu_out_4_ ),
    .B(eu_mdb_out_4_),
    .S(_01127_),
    .Y(_01136_)
  );
  NAND2X1 _07454_ (
    .A(execution_unit_0.pc_nxt_4_ ),
    .B(_01121_),
    .Y(_01137_)
  );
  OAI21X1 _07455_ (
    .A(_01121_),
    .B(_01136_),
    .C(_01137_),
    .Y(_01057_)
  );
  MUX2X1 _07456_ (
    .A(execution_unit_0.alu_0.alu_out_5_ ),
    .B(eu_mdb_out_5_),
    .S(_01127_),
    .Y(_01138_)
  );
  NAND2X1 _07457_ (
    .A(execution_unit_0.pc_nxt_5_ ),
    .B(_01121_),
    .Y(_01139_)
  );
  OAI21X1 _07458_ (
    .A(_01121_),
    .B(_01138_),
    .C(_01139_),
    .Y(_01058_)
  );
  MUX2X1 _07459_ (
    .A(execution_unit_0.alu_0.alu_out_6_ ),
    .B(eu_mdb_out_6_),
    .S(_01127_),
    .Y(_01140_)
  );
  NAND2X1 _07460_ (
    .A(execution_unit_0.pc_nxt_6_ ),
    .B(_01121_),
    .Y(_01141_)
  );
  OAI21X1 _07461_ (
    .A(_01121_),
    .B(_01140_),
    .C(_01141_),
    .Y(_01059_)
  );
  MUX2X1 _07462_ (
    .A(execution_unit_0.alu_0.alu_out_7_ ),
    .B(eu_mdb_out_7_),
    .S(_01127_),
    .Y(_01142_)
  );
  NAND2X1 _07463_ (
    .A(execution_unit_0.pc_nxt_7_ ),
    .B(_01121_),
    .Y(_01143_)
  );
  OAI21X1 _07464_ (
    .A(_01121_),
    .B(_01142_),
    .C(_01143_),
    .Y(_01060_)
  );
  MUX2X1 _07465_ (
    .A(execution_unit_0.alu_0.alu_out_8_ ),
    .B(execution_unit_0.mdb_out_nxt_8_ ),
    .S(_01127_),
    .Y(_01144_)
  );
  NAND2X1 _07466_ (
    .A(execution_unit_0.pc_nxt_8_ ),
    .B(_01121_),
    .Y(_01145_)
  );
  OAI21X1 _07467_ (
    .A(_01121_),
    .B(_01144_),
    .C(_01145_),
    .Y(_01061_)
  );
  MUX2X1 _07468_ (
    .A(execution_unit_0.alu_0.alu_out_9_ ),
    .B(execution_unit_0.mdb_out_nxt_9_ ),
    .S(_01127_),
    .Y(_01146_)
  );
  NAND2X1 _07469_ (
    .A(execution_unit_0.pc_nxt_9_ ),
    .B(_01121_),
    .Y(_01147_)
  );
  OAI21X1 _07470_ (
    .A(_01121_),
    .B(_01146_),
    .C(_01147_),
    .Y(_01062_)
  );
  MUX2X1 _07471_ (
    .A(execution_unit_0.alu_0.alu_out_10_ ),
    .B(execution_unit_0.mdb_out_nxt_10_ ),
    .S(_01127_),
    .Y(_01148_)
  );
  NAND2X1 _07472_ (
    .A(execution_unit_0.pc_nxt_10_ ),
    .B(_01121_),
    .Y(_01149_)
  );
  OAI21X1 _07473_ (
    .A(_01121_),
    .B(_01148_),
    .C(_01149_),
    .Y(_01048_)
  );
  MUX2X1 _07474_ (
    .A(execution_unit_0.alu_0.alu_out_11_ ),
    .B(execution_unit_0.mdb_out_nxt_11_ ),
    .S(_01127_),
    .Y(_01150_)
  );
  NAND2X1 _07475_ (
    .A(execution_unit_0.pc_nxt_11_ ),
    .B(_01121_),
    .Y(_01151_)
  );
  OAI21X1 _07476_ (
    .A(_01121_),
    .B(_01150_),
    .C(_01151_),
    .Y(_01049_)
  );
  MUX2X1 _07477_ (
    .A(execution_unit_0.alu_0.alu_out_12_ ),
    .B(execution_unit_0.mdb_out_nxt_12_ ),
    .S(_01127_),
    .Y(_01152_)
  );
  NAND2X1 _07478_ (
    .A(execution_unit_0.pc_nxt_12_ ),
    .B(_01121_),
    .Y(_01153_)
  );
  OAI21X1 _07479_ (
    .A(_01121_),
    .B(_01152_),
    .C(_01153_),
    .Y(_01050_)
  );
  MUX2X1 _07480_ (
    .A(execution_unit_0.alu_0.alu_out_13_ ),
    .B(execution_unit_0.mdb_out_nxt_13_ ),
    .S(_01127_),
    .Y(_01154_)
  );
  NAND2X1 _07481_ (
    .A(execution_unit_0.pc_nxt_13_ ),
    .B(_01121_),
    .Y(_01155_)
  );
  OAI21X1 _07482_ (
    .A(_01121_),
    .B(_01154_),
    .C(_01155_),
    .Y(_01051_)
  );
  MUX2X1 _07483_ (
    .A(execution_unit_0.alu_0.alu_out_14_ ),
    .B(execution_unit_0.mdb_out_nxt_14_ ),
    .S(_01127_),
    .Y(_01156_)
  );
  NAND2X1 _07484_ (
    .A(execution_unit_0.pc_nxt_14_ ),
    .B(_01121_),
    .Y(_01157_)
  );
  OAI21X1 _07485_ (
    .A(_01121_),
    .B(_01156_),
    .C(_01157_),
    .Y(_01052_)
  );
  MUX2X1 _07486_ (
    .A(execution_unit_0.alu_0.alu_out_15_ ),
    .B(execution_unit_0.mdb_out_nxt_15_ ),
    .S(_01127_),
    .Y(_01158_)
  );
  NAND2X1 _07487_ (
    .A(execution_unit_0.pc_nxt_15_ ),
    .B(_01121_),
    .Y(_01159_)
  );
  OAI21X1 _07488_ (
    .A(_01121_),
    .B(_01158_),
    .C(_01159_),
    .Y(_01053_)
  );
  NOR2X1 _07489_ (
    .A(_01066_),
    .B(_01122_),
    .Y(execution_unit_0.reg_sr_wr )
  );
  NOR2X1 _07490_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B(execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .Y(_01160_)
  );
  OR2X1 _07491_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B(execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .Y(_01161_)
  );
  NOR3X1 _07492_ (
    .A(_01064_),
    .B(e_state_1_),
    .C(_01160_),
    .Y(_01162_)
  );
  NAND2X1 _07493_ (
    .A(_01104_),
    .B(_01162_),
    .Y(_01163_)
  );
  NAND3X1 _07494_ (
    .A(execution_unit_0.inst_as_1_ ),
    .B(_01107_),
    .C(_01162_),
    .Y(_01164_)
  );
  OAI21X1 _07495_ (
    .A(_01122_),
    .B(_01160_),
    .C(_01164_),
    .Y(_01165_)
  );
  AOI21X1 _07496_ (
    .A(e_state_0_),
    .B(_01111_),
    .C(_01165_),
    .Y(_01166_)
  );
  NOR2X1 _07497_ (
    .A(execution_unit_0.inst_as_3_ ),
    .B(execution_unit_0.inst_as_2_ ),
    .Y(_01167_)
  );
  OR2X1 _07498_ (
    .A(execution_unit_0.inst_as_6_ ),
    .B(execution_unit_0.inst_as_1_ ),
    .Y(_01168_)
  );
  NOR2X1 _07499_ (
    .A(execution_unit_0.inst_as_4_ ),
    .B(_01168_),
    .Y(_01169_)
  );
  AOI21X1 _07500_ (
    .A(_01167_),
    .B(_01169_),
    .C(_01106_),
    .Y(_01170_)
  );
  NOR2X1 _07501_ (
    .A(execution_unit_0.reg_sr_wr ),
    .B(_01170_),
    .Y(_01171_)
  );
  AOI21X1 _07502_ (
    .A(_01117_),
    .B(_01122_),
    .C(_01161_),
    .Y(_01172_)
  );
  NOR2X1 _07503_ (
    .A(execution_unit_0.inst_type_1_ ),
    .B(execution_unit_0.inst_as_7_ ),
    .Y(_01173_)
  );
  NOR2X1 _07504_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(execution_unit_0.inst_as_5_ ),
    .Y(_01174_)
  );
  AOI21X1 _07505_ (
    .A(_01173_),
    .B(_01174_),
    .C(_01106_),
    .Y(_01175_)
  );
  AOI22X1 _07506_ (
    .A(execution_unit_0.inst_dext_0_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_0_ ),
    .Y(_01176_)
  );
  NAND2X1 _07507_ (
    .A(execution_unit_0.mab_lsb ),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01177_)
  );
  MUX2X1 _07508_ (
    .A(eu_mdb_in_0_),
    .B(eu_mdb_in_8_),
    .S(_01177_),
    .Y(_01178_)
  );
  NOR2X1 _07509_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01178_),
    .Y(_01179_)
  );
  AOI21X1 _07510_ (
    .A(execution_unit_0.mdb_in_buf_0_ ),
    .B(execution_unit_0.mdb_in_buf_valid ),
    .C(_01179_),
    .Y(_01180_)
  );
  MUX2X1 _07511_ (
    .A(_01176_),
    .B(_01180_),
    .S(_01171_),
    .Y(_01181_)
  );
  NOR2X1 _07512_ (
    .A(execution_unit_0.inst_type_1_ ),
    .B(_01106_),
    .Y(_01182_)
  );
  AOI22X1 _07513_ (
    .A(_01064_),
    .B(_01111_),
    .C(_01182_),
    .D(execution_unit_0.inst_as_0_ ),
    .Y(_01183_)
  );
  OAI21X1 _07514_ (
    .A(execution_unit_0.inst_as_6_ ),
    .B(_01108_),
    .C(_01183_),
    .Y(_01184_)
  );
  MUX2X1 _07515_ (
    .A(_01181_),
    .B(dbg_0.dbg_reg_din_0_ ),
    .S(_01166_),
    .Y(_01185_)
  );
  NAND2X1 _07516_ (
    .A(execution_unit_0.reg_src_0_ ),
    .B(_01184_),
    .Y(_01186_)
  );
  OAI21X1 _07517_ (
    .A(_01184_),
    .B(_01185_),
    .C(_01186_),
    .Y(execution_unit_0.alu_0.alu_swpb_8_ )
  );
  AOI22X1 _07518_ (
    .A(execution_unit_0.inst_dext_1_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_1_ ),
    .Y(_01187_)
  );
  MUX2X1 _07519_ (
    .A(eu_mdb_in_1_),
    .B(eu_mdb_in_9_),
    .S(_01177_),
    .Y(_01188_)
  );
  NOR2X1 _07520_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01188_),
    .Y(_01189_)
  );
  AOI21X1 _07521_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(execution_unit_0.mdb_in_buf_1_ ),
    .C(_01189_),
    .Y(_01190_)
  );
  MUX2X1 _07522_ (
    .A(_01187_),
    .B(_01190_),
    .S(_01171_),
    .Y(_01191_)
  );
  MUX2X1 _07523_ (
    .A(_01191_),
    .B(dbg_0.dbg_reg_din_1_ ),
    .S(_01166_),
    .Y(_01192_)
  );
  NAND2X1 _07524_ (
    .A(execution_unit_0.reg_src_1_ ),
    .B(_01184_),
    .Y(_01193_)
  );
  OAI21X1 _07525_ (
    .A(_01184_),
    .B(_01192_),
    .C(_01193_),
    .Y(execution_unit_0.alu_0.alu_shift_0_ )
  );
  AOI22X1 _07526_ (
    .A(execution_unit_0.inst_dext_2_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_2_ ),
    .Y(_01194_)
  );
  MUX2X1 _07527_ (
    .A(eu_mdb_in_2_),
    .B(eu_mdb_in_10_),
    .S(_01177_),
    .Y(_01195_)
  );
  NOR2X1 _07528_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01195_),
    .Y(_01196_)
  );
  AOI21X1 _07529_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(execution_unit_0.mdb_in_buf_2_ ),
    .C(_01196_),
    .Y(_01197_)
  );
  MUX2X1 _07530_ (
    .A(_01194_),
    .B(_01197_),
    .S(_01171_),
    .Y(_01198_)
  );
  MUX2X1 _07531_ (
    .A(_01198_),
    .B(dbg_0.dbg_reg_din_2_ ),
    .S(_01166_),
    .Y(_01199_)
  );
  NAND2X1 _07532_ (
    .A(execution_unit_0.reg_src_2_ ),
    .B(_01184_),
    .Y(_01200_)
  );
  OAI21X1 _07533_ (
    .A(_01184_),
    .B(_01199_),
    .C(_01200_),
    .Y(execution_unit_0.alu_0.alu_shift_1_ )
  );
  AOI22X1 _07534_ (
    .A(execution_unit_0.inst_dext_3_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_3_ ),
    .Y(_01201_)
  );
  MUX2X1 _07535_ (
    .A(eu_mdb_in_3_),
    .B(eu_mdb_in_11_),
    .S(_01177_),
    .Y(_01202_)
  );
  NOR2X1 _07536_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01202_),
    .Y(_01203_)
  );
  AOI21X1 _07537_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(execution_unit_0.mdb_in_buf_3_ ),
    .C(_01203_),
    .Y(_01204_)
  );
  MUX2X1 _07538_ (
    .A(_01201_),
    .B(_01204_),
    .S(_01171_),
    .Y(_01205_)
  );
  MUX2X1 _07539_ (
    .A(_01205_),
    .B(dbg_0.dbg_reg_din_3_ ),
    .S(_01166_),
    .Y(_01206_)
  );
  NAND2X1 _07540_ (
    .A(execution_unit_0.reg_src_3_ ),
    .B(_01184_),
    .Y(_01207_)
  );
  OAI21X1 _07541_ (
    .A(_01184_),
    .B(_01206_),
    .C(_01207_),
    .Y(execution_unit_0.alu_0.alu_shift_2_ )
  );
  AOI22X1 _07542_ (
    .A(execution_unit_0.inst_dext_4_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_4_ ),
    .Y(_01208_)
  );
  MUX2X1 _07543_ (
    .A(eu_mdb_in_4_),
    .B(eu_mdb_in_12_),
    .S(_01177_),
    .Y(_01209_)
  );
  NOR2X1 _07544_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01209_),
    .Y(_01210_)
  );
  AOI21X1 _07545_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(execution_unit_0.mdb_in_buf_4_ ),
    .C(_01210_),
    .Y(_01211_)
  );
  MUX2X1 _07546_ (
    .A(_01208_),
    .B(_01211_),
    .S(_01171_),
    .Y(_01212_)
  );
  MUX2X1 _07547_ (
    .A(_01212_),
    .B(dbg_0.dbg_reg_din_4_ ),
    .S(_01166_),
    .Y(_01213_)
  );
  NAND2X1 _07548_ (
    .A(execution_unit_0.reg_src_4_ ),
    .B(_01184_),
    .Y(_01214_)
  );
  OAI21X1 _07549_ (
    .A(_01184_),
    .B(_01213_),
    .C(_01214_),
    .Y(execution_unit_0.alu_0.alu_shift_3_ )
  );
  AOI22X1 _07550_ (
    .A(execution_unit_0.inst_dext_5_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_5_ ),
    .Y(_01215_)
  );
  MUX2X1 _07551_ (
    .A(eu_mdb_in_5_),
    .B(eu_mdb_in_13_),
    .S(_01177_),
    .Y(_01216_)
  );
  NOR2X1 _07552_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01216_),
    .Y(_01217_)
  );
  AOI21X1 _07553_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(execution_unit_0.mdb_in_buf_5_ ),
    .C(_01217_),
    .Y(_01218_)
  );
  MUX2X1 _07554_ (
    .A(_01215_),
    .B(_01218_),
    .S(_01171_),
    .Y(_01219_)
  );
  MUX2X1 _07555_ (
    .A(_01219_),
    .B(dbg_0.dbg_reg_din_5_ ),
    .S(_01166_),
    .Y(_01220_)
  );
  NAND2X1 _07556_ (
    .A(execution_unit_0.reg_src_5_ ),
    .B(_01184_),
    .Y(_01221_)
  );
  OAI21X1 _07557_ (
    .A(_01184_),
    .B(_01220_),
    .C(_01221_),
    .Y(execution_unit_0.alu_0.alu_shift_4_ )
  );
  AOI22X1 _07558_ (
    .A(execution_unit_0.inst_dext_6_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_6_ ),
    .Y(_01222_)
  );
  MUX2X1 _07559_ (
    .A(eu_mdb_in_6_),
    .B(eu_mdb_in_14_),
    .S(_01177_),
    .Y(_01223_)
  );
  NOR2X1 _07560_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01223_),
    .Y(_01224_)
  );
  AOI21X1 _07561_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(execution_unit_0.mdb_in_buf_6_ ),
    .C(_01224_),
    .Y(_01225_)
  );
  MUX2X1 _07562_ (
    .A(_01222_),
    .B(_01225_),
    .S(_01171_),
    .Y(_01226_)
  );
  MUX2X1 _07563_ (
    .A(_01226_),
    .B(dbg_0.dbg_reg_din_6_ ),
    .S(_01166_),
    .Y(_01227_)
  );
  NAND2X1 _07564_ (
    .A(execution_unit_0.reg_src_6_ ),
    .B(_01184_),
    .Y(_01228_)
  );
  OAI21X1 _07565_ (
    .A(_01184_),
    .B(_01227_),
    .C(_01228_),
    .Y(execution_unit_0.alu_0.alu_shift_5_ )
  );
  AOI22X1 _07566_ (
    .A(execution_unit_0.inst_dext_7_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_7_ ),
    .Y(_01229_)
  );
  MUX2X1 _07567_ (
    .A(eu_mdb_in_7_),
    .B(eu_mdb_in_15_),
    .S(_01177_),
    .Y(_01230_)
  );
  NOR2X1 _07568_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01230_),
    .Y(_01231_)
  );
  AOI21X1 _07569_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(execution_unit_0.mdb_in_buf_7_ ),
    .C(_01231_),
    .Y(_01232_)
  );
  MUX2X1 _07570_ (
    .A(_01229_),
    .B(_01232_),
    .S(_01171_),
    .Y(_01233_)
  );
  MUX2X1 _07571_ (
    .A(_01233_),
    .B(dbg_0.dbg_reg_din_7_ ),
    .S(_01166_),
    .Y(_01234_)
  );
  NAND2X1 _07572_ (
    .A(execution_unit_0.reg_src_7_ ),
    .B(_01184_),
    .Y(_01235_)
  );
  OAI21X1 _07573_ (
    .A(_01184_),
    .B(_01234_),
    .C(_01235_),
    .Y(execution_unit_0.alu_0.alu_shift_6_ )
  );
  AOI22X1 _07574_ (
    .A(execution_unit_0.inst_dext_8_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_8_ ),
    .Y(_01236_)
  );
  MUX2X1 _07575_ (
    .A(execution_unit_0.mdb_in_buf_8_ ),
    .B(eu_mdb_in_8_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01237_)
  );
  MUX2X1 _07576_ (
    .A(_01236_),
    .B(_01237_),
    .S(_01171_),
    .Y(_01238_)
  );
  MUX2X1 _07577_ (
    .A(_01238_),
    .B(dbg_0.dbg_reg_din_8_ ),
    .S(_01166_),
    .Y(_01239_)
  );
  NAND2X1 _07578_ (
    .A(execution_unit_0.reg_src_8_ ),
    .B(_01184_),
    .Y(_01240_)
  );
  OAI21X1 _07579_ (
    .A(_01184_),
    .B(_01239_),
    .C(_01240_),
    .Y(execution_unit_0.alu_0.alu_swpb_0_ )
  );
  AOI22X1 _07580_ (
    .A(execution_unit_0.inst_dext_9_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_9_ ),
    .Y(_01241_)
  );
  MUX2X1 _07581_ (
    .A(execution_unit_0.mdb_in_buf_9_ ),
    .B(eu_mdb_in_9_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01242_)
  );
  MUX2X1 _07582_ (
    .A(_01241_),
    .B(_01242_),
    .S(_01171_),
    .Y(_01243_)
  );
  MUX2X1 _07583_ (
    .A(_01243_),
    .B(dbg_0.dbg_reg_din_9_ ),
    .S(_01166_),
    .Y(_01244_)
  );
  NAND2X1 _07584_ (
    .A(execution_unit_0.reg_src_9_ ),
    .B(_01184_),
    .Y(_01245_)
  );
  OAI21X1 _07585_ (
    .A(_01184_),
    .B(_01244_),
    .C(_01245_),
    .Y(execution_unit_0.alu_0.alu_shift_8_ )
  );
  AOI22X1 _07586_ (
    .A(execution_unit_0.inst_dext_10_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_10_ ),
    .Y(_01246_)
  );
  MUX2X1 _07587_ (
    .A(execution_unit_0.mdb_in_buf_10_ ),
    .B(eu_mdb_in_10_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01247_)
  );
  MUX2X1 _07588_ (
    .A(_01246_),
    .B(_01247_),
    .S(_01171_),
    .Y(_01248_)
  );
  MUX2X1 _07589_ (
    .A(_01248_),
    .B(dbg_0.dbg_reg_din_10_ ),
    .S(_01166_),
    .Y(_01249_)
  );
  NAND2X1 _07590_ (
    .A(execution_unit_0.reg_src_10_ ),
    .B(_01184_),
    .Y(_01250_)
  );
  OAI21X1 _07591_ (
    .A(_01184_),
    .B(_01249_),
    .C(_01250_),
    .Y(execution_unit_0.alu_0.alu_shift_9_ )
  );
  AOI22X1 _07592_ (
    .A(execution_unit_0.inst_dext_11_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_11_ ),
    .Y(_01251_)
  );
  MUX2X1 _07593_ (
    .A(execution_unit_0.mdb_in_buf_11_ ),
    .B(eu_mdb_in_11_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01252_)
  );
  MUX2X1 _07594_ (
    .A(_01251_),
    .B(_01252_),
    .S(_01171_),
    .Y(_01253_)
  );
  MUX2X1 _07595_ (
    .A(_01253_),
    .B(dbg_0.dbg_reg_din_11_ ),
    .S(_01166_),
    .Y(_01254_)
  );
  NAND2X1 _07596_ (
    .A(execution_unit_0.reg_src_11_ ),
    .B(_01184_),
    .Y(_01255_)
  );
  OAI21X1 _07597_ (
    .A(_01184_),
    .B(_01254_),
    .C(_01255_),
    .Y(execution_unit_0.alu_0.alu_shift_10_ )
  );
  AOI22X1 _07598_ (
    .A(execution_unit_0.inst_dext_12_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_12_ ),
    .Y(_01256_)
  );
  MUX2X1 _07599_ (
    .A(execution_unit_0.mdb_in_buf_12_ ),
    .B(eu_mdb_in_12_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01257_)
  );
  MUX2X1 _07600_ (
    .A(_01256_),
    .B(_01257_),
    .S(_01171_),
    .Y(_01258_)
  );
  MUX2X1 _07601_ (
    .A(_01258_),
    .B(dbg_0.dbg_reg_din_12_ ),
    .S(_01166_),
    .Y(_01259_)
  );
  NAND2X1 _07602_ (
    .A(execution_unit_0.reg_src_12_ ),
    .B(_01184_),
    .Y(_01260_)
  );
  OAI21X1 _07603_ (
    .A(_01184_),
    .B(_01259_),
    .C(_01260_),
    .Y(execution_unit_0.alu_0.alu_shift_11_ )
  );
  AOI22X1 _07604_ (
    .A(execution_unit_0.inst_dext_13_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_13_ ),
    .Y(_01261_)
  );
  MUX2X1 _07605_ (
    .A(execution_unit_0.mdb_in_buf_13_ ),
    .B(eu_mdb_in_13_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01262_)
  );
  MUX2X1 _07606_ (
    .A(_01261_),
    .B(_01262_),
    .S(_01171_),
    .Y(_01263_)
  );
  MUX2X1 _07607_ (
    .A(_01263_),
    .B(dbg_0.dbg_reg_din_13_ ),
    .S(_01166_),
    .Y(_01264_)
  );
  NAND2X1 _07608_ (
    .A(execution_unit_0.reg_src_13_ ),
    .B(_01184_),
    .Y(_01265_)
  );
  OAI21X1 _07609_ (
    .A(_01184_),
    .B(_01264_),
    .C(_01265_),
    .Y(execution_unit_0.alu_0.alu_shift_12_ )
  );
  AOI22X1 _07610_ (
    .A(execution_unit_0.inst_dext_14_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_14_ ),
    .Y(_01266_)
  );
  MUX2X1 _07611_ (
    .A(execution_unit_0.mdb_in_buf_14_ ),
    .B(eu_mdb_in_14_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01267_)
  );
  MUX2X1 _07612_ (
    .A(_01266_),
    .B(_01267_),
    .S(_01171_),
    .Y(_01268_)
  );
  MUX2X1 _07613_ (
    .A(_01268_),
    .B(dbg_0.dbg_reg_din_14_ ),
    .S(_01166_),
    .Y(_01269_)
  );
  NAND2X1 _07614_ (
    .A(execution_unit_0.reg_src_14_ ),
    .B(_01184_),
    .Y(_01270_)
  );
  OAI21X1 _07615_ (
    .A(_01184_),
    .B(_01269_),
    .C(_01270_),
    .Y(execution_unit_0.alu_0.alu_shift_13_ )
  );
  AOI22X1 _07616_ (
    .A(execution_unit_0.inst_dext_15_ ),
    .B(_01172_),
    .C(_01175_),
    .D(execution_unit_0.inst_sext_15_ ),
    .Y(_01271_)
  );
  MUX2X1 _07617_ (
    .A(execution_unit_0.mdb_in_buf_15_ ),
    .B(eu_mdb_in_15_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01272_)
  );
  MUX2X1 _07618_ (
    .A(_01271_),
    .B(_01272_),
    .S(_01171_),
    .Y(_01273_)
  );
  MUX2X1 _07619_ (
    .A(_01273_),
    .B(dbg_0.dbg_reg_din_15_ ),
    .S(_01166_),
    .Y(_01274_)
  );
  NAND2X1 _07620_ (
    .A(execution_unit_0.reg_src_15_ ),
    .B(_01184_),
    .Y(_01275_)
  );
  OAI21X1 _07621_ (
    .A(_01184_),
    .B(_01274_),
    .C(_01275_),
    .Y(execution_unit_0.alu_0.alu_shift_14_ )
  );
  OR2X1 _07622_ (
    .A(execution_unit_0.inst_type_0_ ),
    .B(execution_unit_0.inst_type_1_ ),
    .Y(_01276_)
  );
  NOR2X1 _07623_ (
    .A(execution_unit_0.inst_ad_0_ ),
    .B(_01276_),
    .Y(_01277_)
  );
  INVX1 _07624_ (
    .A(_01277_),
    .Y(_01278_)
  );
  OR2X1 _07625_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01106_),
    .Y(_01279_)
  );
  NOR2X1 _07626_ (
    .A(_01277_),
    .B(_01279_),
    .Y(_01280_)
  );
  NOR2X1 _07627_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01161_),
    .Y(_01281_)
  );
  NAND3X1 _07628_ (
    .A(_01104_),
    .B(_01120_),
    .C(_01281_),
    .Y(_01282_)
  );
  AOI21X1 _07629_ (
    .A(_01116_),
    .B(_01282_),
    .C(execution_unit_0.inst_ad_6_ ),
    .Y(_01283_)
  );
  NOR2X1 _07630_ (
    .A(_01280_),
    .B(_01283_),
    .Y(_01284_)
  );
  NOR2X1 _07631_ (
    .A(_01278_),
    .B(_01279_),
    .Y(_01285_)
  );
  NAND3X1 _07632_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01104_),
    .C(_01109_),
    .Y(_01286_)
  );
  INVX1 _07633_ (
    .A(_01286_),
    .Y(_01287_)
  );
  NOR2X1 _07634_ (
    .A(_01285_),
    .B(_01287_),
    .Y(_01288_)
  );
  OAI21X1 _07635_ (
    .A(_01278_),
    .B(_01279_),
    .C(_01286_),
    .Y(_01289_)
  );
  NOR2X1 _07636_ (
    .A(_01284_),
    .B(_01289_),
    .Y(_01290_)
  );
  NOR2X1 _07637_ (
    .A(_01108_),
    .B(_01169_),
    .Y(_01291_)
  );
  OR2X1 _07638_ (
    .A(_01108_),
    .B(_01169_),
    .Y(_01292_)
  );
  NAND2X1 _07639_ (
    .A(execution_unit_0.inst_sext_0_ ),
    .B(_01291_),
    .Y(_01293_)
  );
  OAI21X1 _07640_ (
    .A(_01178_),
    .B(_01288_),
    .C(_01293_),
    .Y(_01294_)
  );
  AOI21X1 _07641_ (
    .A(dbg_0.dbg_reg_din_0_ ),
    .B(_01290_),
    .C(_01294_),
    .Y(_01295_)
  );
  NAND2X1 _07642_ (
    .A(_00144_),
    .B(cpu_halt_st),
    .Y(_01296_)
  );
  OAI21X1 _07643_ (
    .A(cpu_halt_st),
    .B(_01295_),
    .C(_01296_),
    .Y(execution_unit_0.alu_0.op_dst_0_ )
  );
  NAND2X1 _07644_ (
    .A(cpu_halt_st),
    .B(_00151_),
    .Y(_01297_)
  );
  OAI21X1 _07645_ (
    .A(execution_unit_0.inst_as_3_ ),
    .B(execution_unit_0.inst_as_2_ ),
    .C(execution_unit_0.inst_src_1_ ),
    .Y(_01298_)
  );
  INVX1 _07646_ (
    .A(_01298_),
    .Y(_01299_)
  );
  OAI21X1 _07647_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B(execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .C(_01299_),
    .Y(_01300_)
  );
  OAI21X1 _07648_ (
    .A(_01110_),
    .B(_01300_),
    .C(_01164_),
    .Y(_01301_)
  );
  OAI21X1 _07649_ (
    .A(e_state_0_),
    .B(e_state_1_),
    .C(_01111_),
    .Y(_01302_)
  );
  OAI21X1 _07650_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01163_),
    .C(_01302_),
    .Y(_01303_)
  );
  NOR3X1 _07651_ (
    .A(_01289_),
    .B(_01301_),
    .C(_01303_),
    .Y(_01304_)
  );
  OAI21X1 _07652_ (
    .A(_01079_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01305_)
  );
  OAI21X1 _07653_ (
    .A(_01285_),
    .B(_01287_),
    .C(_01188_),
    .Y(_01306_)
  );
  AOI21X1 _07654_ (
    .A(_01305_),
    .B(_01306_),
    .C(_01291_),
    .Y(_01307_)
  );
  OAI21X1 _07655_ (
    .A(execution_unit_0.inst_sext_1_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01308_)
  );
  OAI21X1 _07656_ (
    .A(_01307_),
    .B(_01308_),
    .C(_01297_),
    .Y(execution_unit_0.alu_0.op_dst_1_ )
  );
  NAND2X1 _07657_ (
    .A(cpu_halt_st),
    .B(_00152_),
    .Y(_01309_)
  );
  OAI21X1 _07658_ (
    .A(_01080_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01310_)
  );
  OAI21X1 _07659_ (
    .A(_01285_),
    .B(_01287_),
    .C(_01195_),
    .Y(_01311_)
  );
  AOI21X1 _07660_ (
    .A(_01310_),
    .B(_01311_),
    .C(_01291_),
    .Y(_01312_)
  );
  OAI21X1 _07661_ (
    .A(execution_unit_0.inst_sext_2_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01313_)
  );
  OAI21X1 _07662_ (
    .A(_01312_),
    .B(_01313_),
    .C(_01309_),
    .Y(execution_unit_0.alu_0.op_dst_2_ )
  );
  NAND2X1 _07663_ (
    .A(cpu_halt_st),
    .B(_00153_),
    .Y(_01314_)
  );
  OAI21X1 _07664_ (
    .A(_01081_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01315_)
  );
  OAI21X1 _07665_ (
    .A(_01285_),
    .B(_01287_),
    .C(_01202_),
    .Y(_01316_)
  );
  AOI21X1 _07666_ (
    .A(_01315_),
    .B(_01316_),
    .C(_01291_),
    .Y(_01317_)
  );
  OAI21X1 _07667_ (
    .A(execution_unit_0.inst_sext_3_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01318_)
  );
  OAI21X1 _07668_ (
    .A(_01317_),
    .B(_01318_),
    .C(_01314_),
    .Y(execution_unit_0.alu_0.op_dst_3_ )
  );
  NAND2X1 _07669_ (
    .A(cpu_halt_st),
    .B(_00154_),
    .Y(_01319_)
  );
  OAI21X1 _07670_ (
    .A(_01082_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01320_)
  );
  OAI21X1 _07671_ (
    .A(_01285_),
    .B(_01287_),
    .C(_01209_),
    .Y(_01321_)
  );
  AOI21X1 _07672_ (
    .A(_01320_),
    .B(_01321_),
    .C(_01291_),
    .Y(_01322_)
  );
  OAI21X1 _07673_ (
    .A(execution_unit_0.inst_sext_4_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01323_)
  );
  OAI21X1 _07674_ (
    .A(_01322_),
    .B(_01323_),
    .C(_01319_),
    .Y(execution_unit_0.alu_0.op_dst_4_ )
  );
  NAND2X1 _07675_ (
    .A(cpu_halt_st),
    .B(_00155_),
    .Y(_01324_)
  );
  OAI21X1 _07676_ (
    .A(_01083_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01325_)
  );
  OAI21X1 _07677_ (
    .A(_01285_),
    .B(_01287_),
    .C(_01216_),
    .Y(_01326_)
  );
  AOI21X1 _07678_ (
    .A(_01325_),
    .B(_01326_),
    .C(_01291_),
    .Y(_01327_)
  );
  OAI21X1 _07679_ (
    .A(execution_unit_0.inst_sext_5_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01328_)
  );
  OAI21X1 _07680_ (
    .A(_01327_),
    .B(_01328_),
    .C(_01324_),
    .Y(execution_unit_0.alu_0.op_dst_5_ )
  );
  NAND2X1 _07681_ (
    .A(cpu_halt_st),
    .B(_00156_),
    .Y(_01329_)
  );
  OAI21X1 _07682_ (
    .A(_01084_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01330_)
  );
  OAI21X1 _07683_ (
    .A(_01285_),
    .B(_01287_),
    .C(_01223_),
    .Y(_01331_)
  );
  AOI21X1 _07684_ (
    .A(_01330_),
    .B(_01331_),
    .C(_01291_),
    .Y(_01332_)
  );
  OAI21X1 _07685_ (
    .A(execution_unit_0.inst_sext_6_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01333_)
  );
  OAI21X1 _07686_ (
    .A(_01332_),
    .B(_01333_),
    .C(_01329_),
    .Y(execution_unit_0.alu_0.op_dst_6_ )
  );
  NAND2X1 _07687_ (
    .A(cpu_halt_st),
    .B(_00157_),
    .Y(_01334_)
  );
  OAI21X1 _07688_ (
    .A(_01085_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01335_)
  );
  OAI21X1 _07689_ (
    .A(_01285_),
    .B(_01287_),
    .C(_01230_),
    .Y(_01336_)
  );
  AOI21X1 _07690_ (
    .A(_01335_),
    .B(_01336_),
    .C(_01291_),
    .Y(_01337_)
  );
  OAI21X1 _07691_ (
    .A(execution_unit_0.inst_sext_7_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01338_)
  );
  OAI21X1 _07692_ (
    .A(_01337_),
    .B(_01338_),
    .C(_01334_),
    .Y(execution_unit_0.alu_0.op_dst_7_ )
  );
  NAND2X1 _07693_ (
    .A(cpu_halt_st),
    .B(_00158_),
    .Y(_01339_)
  );
  OAI21X1 _07694_ (
    .A(_01087_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01340_)
  );
  OR2X1 _07695_ (
    .A(eu_mdb_in_8_),
    .B(_01288_),
    .Y(_01341_)
  );
  AOI21X1 _07696_ (
    .A(_01340_),
    .B(_01341_),
    .C(_01291_),
    .Y(_01342_)
  );
  OAI21X1 _07697_ (
    .A(execution_unit_0.inst_sext_8_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01343_)
  );
  OAI21X1 _07698_ (
    .A(_01342_),
    .B(_01343_),
    .C(_01339_),
    .Y(execution_unit_0.alu_0.op_dst_8_ )
  );
  NAND2X1 _07699_ (
    .A(cpu_halt_st),
    .B(_00159_),
    .Y(_01344_)
  );
  OAI21X1 _07700_ (
    .A(_01089_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01345_)
  );
  OR2X1 _07701_ (
    .A(eu_mdb_in_9_),
    .B(_01288_),
    .Y(_01346_)
  );
  AOI21X1 _07702_ (
    .A(_01345_),
    .B(_01346_),
    .C(_01291_),
    .Y(_01347_)
  );
  OAI21X1 _07703_ (
    .A(execution_unit_0.inst_sext_9_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01348_)
  );
  OAI21X1 _07704_ (
    .A(_01347_),
    .B(_01348_),
    .C(_01344_),
    .Y(execution_unit_0.alu_0.op_dst_9_ )
  );
  NAND2X1 _07705_ (
    .A(cpu_halt_st),
    .B(_00145_),
    .Y(_01349_)
  );
  OAI21X1 _07706_ (
    .A(_01091_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01350_)
  );
  OR2X1 _07707_ (
    .A(eu_mdb_in_10_),
    .B(_01288_),
    .Y(_01351_)
  );
  AOI21X1 _07708_ (
    .A(_01350_),
    .B(_01351_),
    .C(_01291_),
    .Y(_01352_)
  );
  OAI21X1 _07709_ (
    .A(execution_unit_0.inst_sext_10_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01353_)
  );
  OAI21X1 _07710_ (
    .A(_01352_),
    .B(_01353_),
    .C(_01349_),
    .Y(execution_unit_0.alu_0.op_dst_10_ )
  );
  NAND2X1 _07711_ (
    .A(cpu_halt_st),
    .B(_00146_),
    .Y(_01354_)
  );
  OAI21X1 _07712_ (
    .A(_01093_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01355_)
  );
  OR2X1 _07713_ (
    .A(eu_mdb_in_11_),
    .B(_01288_),
    .Y(_01356_)
  );
  AOI21X1 _07714_ (
    .A(_01355_),
    .B(_01356_),
    .C(_01291_),
    .Y(_01357_)
  );
  OAI21X1 _07715_ (
    .A(execution_unit_0.inst_sext_11_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01358_)
  );
  OAI21X1 _07716_ (
    .A(_01357_),
    .B(_01358_),
    .C(_01354_),
    .Y(execution_unit_0.alu_0.op_dst_11_ )
  );
  NAND2X1 _07717_ (
    .A(cpu_halt_st),
    .B(_00147_),
    .Y(_01359_)
  );
  OAI21X1 _07718_ (
    .A(_01095_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01360_)
  );
  OR2X1 _07719_ (
    .A(eu_mdb_in_12_),
    .B(_01288_),
    .Y(_01361_)
  );
  AOI21X1 _07720_ (
    .A(_01360_),
    .B(_01361_),
    .C(_01291_),
    .Y(_01362_)
  );
  OAI21X1 _07721_ (
    .A(execution_unit_0.inst_sext_12_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01363_)
  );
  OAI21X1 _07722_ (
    .A(_01362_),
    .B(_01363_),
    .C(_01359_),
    .Y(execution_unit_0.alu_0.op_dst_12_ )
  );
  NAND2X1 _07723_ (
    .A(cpu_halt_st),
    .B(_00148_),
    .Y(_01364_)
  );
  OAI21X1 _07724_ (
    .A(_01097_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01365_)
  );
  OR2X1 _07725_ (
    .A(eu_mdb_in_13_),
    .B(_01288_),
    .Y(_01366_)
  );
  AOI21X1 _07726_ (
    .A(_01365_),
    .B(_01366_),
    .C(_01291_),
    .Y(_01367_)
  );
  OAI21X1 _07727_ (
    .A(execution_unit_0.inst_sext_13_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01368_)
  );
  OAI21X1 _07728_ (
    .A(_01367_),
    .B(_01368_),
    .C(_01364_),
    .Y(execution_unit_0.alu_0.op_dst_13_ )
  );
  NAND2X1 _07729_ (
    .A(cpu_halt_st),
    .B(_00149_),
    .Y(_01369_)
  );
  OAI21X1 _07730_ (
    .A(_01099_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01370_)
  );
  OR2X1 _07731_ (
    .A(eu_mdb_in_14_),
    .B(_01288_),
    .Y(_01371_)
  );
  AOI21X1 _07732_ (
    .A(_01370_),
    .B(_01371_),
    .C(_01291_),
    .Y(_01372_)
  );
  OAI21X1 _07733_ (
    .A(execution_unit_0.inst_sext_14_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01373_)
  );
  OAI21X1 _07734_ (
    .A(_01372_),
    .B(_01373_),
    .C(_01369_),
    .Y(execution_unit_0.alu_0.op_dst_14_ )
  );
  NAND2X1 _07735_ (
    .A(cpu_halt_st),
    .B(_00150_),
    .Y(_01374_)
  );
  OAI21X1 _07736_ (
    .A(_01101_),
    .B(_01284_),
    .C(_01304_),
    .Y(_01375_)
  );
  OR2X1 _07737_ (
    .A(eu_mdb_in_15_),
    .B(_01288_),
    .Y(_01376_)
  );
  AOI21X1 _07738_ (
    .A(_01375_),
    .B(_01376_),
    .C(_01291_),
    .Y(_01377_)
  );
  OAI21X1 _07739_ (
    .A(execution_unit_0.inst_sext_15_ ),
    .B(_01292_),
    .C(_01102_),
    .Y(_01378_)
  );
  OAI21X1 _07740_ (
    .A(_01377_),
    .B(_01378_),
    .C(_01374_),
    .Y(execution_unit_0.alu_0.op_dst_15_ )
  );
  NAND2X1 _07741_ (
    .A(eu_mdb_out_0_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01379_)
  );
  OAI21X1 _07742_ (
    .A(_01071_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01379_),
    .Y(eu_mdb_out_8_)
  );
  NAND2X1 _07743_ (
    .A(eu_mdb_out_1_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01380_)
  );
  OAI21X1 _07744_ (
    .A(_01072_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01380_),
    .Y(eu_mdb_out_9_)
  );
  NAND2X1 _07745_ (
    .A(eu_mdb_out_2_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01381_)
  );
  OAI21X1 _07746_ (
    .A(_01073_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01381_),
    .Y(eu_mdb_out_10_)
  );
  NAND2X1 _07747_ (
    .A(eu_mdb_out_3_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01382_)
  );
  OAI21X1 _07748_ (
    .A(_01074_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01382_),
    .Y(eu_mdb_out_11_)
  );
  NAND2X1 _07749_ (
    .A(eu_mdb_out_4_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01383_)
  );
  OAI21X1 _07750_ (
    .A(_01075_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01383_),
    .Y(eu_mdb_out_12_)
  );
  NAND2X1 _07751_ (
    .A(eu_mdb_out_5_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01384_)
  );
  OAI21X1 _07752_ (
    .A(_01076_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01384_),
    .Y(eu_mdb_out_13_)
  );
  NAND2X1 _07753_ (
    .A(eu_mdb_out_6_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01385_)
  );
  OAI21X1 _07754_ (
    .A(_01077_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01385_),
    .Y(eu_mdb_out_14_)
  );
  NAND2X1 _07755_ (
    .A(eu_mdb_out_7_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01386_)
  );
  OAI21X1 _07756_ (
    .A(_01078_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01386_),
    .Y(eu_mdb_out_15_)
  );
  OAI21X1 _07757_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(execution_unit_0.mdb_in_buf_en ),
    .C(_01106_),
    .Y(_01387_)
  );
  INVX1 _07758_ (
    .A(_01387_),
    .Y(_01046_)
  );
  NOR2X1 _07759_ (
    .A(execution_unit_0.mdb_in_buf_0_ ),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01388_)
  );
  AOI21X1 _07760_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01178_),
    .C(_01388_),
    .Y(_01029_)
  );
  NOR2X1 _07761_ (
    .A(execution_unit_0.mdb_in_buf_1_ ),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01389_)
  );
  AOI21X1 _07762_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01188_),
    .C(_01389_),
    .Y(_01036_)
  );
  NOR2X1 _07763_ (
    .A(execution_unit_0.mdb_in_buf_2_ ),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01390_)
  );
  AOI21X1 _07764_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01195_),
    .C(_01390_),
    .Y(_01037_)
  );
  NOR2X1 _07765_ (
    .A(execution_unit_0.mdb_in_buf_3_ ),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01391_)
  );
  AOI21X1 _07766_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01202_),
    .C(_01391_),
    .Y(_01038_)
  );
  NOR2X1 _07767_ (
    .A(execution_unit_0.mdb_in_buf_4_ ),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01392_)
  );
  AOI21X1 _07768_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01209_),
    .C(_01392_),
    .Y(_01039_)
  );
  NOR2X1 _07769_ (
    .A(execution_unit_0.mdb_in_buf_5_ ),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01393_)
  );
  AOI21X1 _07770_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01216_),
    .C(_01393_),
    .Y(_01040_)
  );
  NOR2X1 _07771_ (
    .A(execution_unit_0.mdb_in_buf_6_ ),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01394_)
  );
  AOI21X1 _07772_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01223_),
    .C(_01394_),
    .Y(_01041_)
  );
  NOR2X1 _07773_ (
    .A(execution_unit_0.mdb_in_buf_7_ ),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01395_)
  );
  AOI21X1 _07774_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01230_),
    .C(_01395_),
    .Y(_01042_)
  );
  NAND2X1 _07775_ (
    .A(eu_mdb_in_8_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01396_)
  );
  OAI21X1 _07776_ (
    .A(_01086_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .C(_01396_),
    .Y(_01043_)
  );
  NAND2X1 _07777_ (
    .A(eu_mdb_in_9_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01397_)
  );
  OAI21X1 _07778_ (
    .A(_01088_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .C(_01397_),
    .Y(_01044_)
  );
  NAND2X1 _07779_ (
    .A(eu_mdb_in_10_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01398_)
  );
  OAI21X1 _07780_ (
    .A(_01090_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .C(_01398_),
    .Y(_01030_)
  );
  NAND2X1 _07781_ (
    .A(eu_mdb_in_11_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01399_)
  );
  OAI21X1 _07782_ (
    .A(_01092_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .C(_01399_),
    .Y(_01031_)
  );
  NAND2X1 _07783_ (
    .A(eu_mdb_in_12_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01400_)
  );
  OAI21X1 _07784_ (
    .A(_01094_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .C(_01400_),
    .Y(_01032_)
  );
  NAND2X1 _07785_ (
    .A(eu_mdb_in_13_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01401_)
  );
  OAI21X1 _07786_ (
    .A(_01096_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .C(_01401_),
    .Y(_01033_)
  );
  NAND2X1 _07787_ (
    .A(eu_mdb_in_14_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01402_)
  );
  OAI21X1 _07788_ (
    .A(_01098_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .C(_01402_),
    .Y(_01034_)
  );
  NAND2X1 _07789_ (
    .A(eu_mdb_in_15_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01403_)
  );
  OAI21X1 _07790_ (
    .A(_01100_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .C(_01403_),
    .Y(_01035_)
  );
  NAND3X1 _07791_ (
    .A(execution_unit_0.inst_type_0_ ),
    .B(execution_unit_0.inst_as_0_ ),
    .C(_01281_),
    .Y(_01404_)
  );
  NAND2X1 _07792_ (
    .A(execution_unit_0.inst_ad_0_ ),
    .B(execution_unit_0.inst_type_2_ ),
    .Y(_01405_)
  );
  OAI21X1 _07793_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_alu ),
    .B(_01405_),
    .C(_01404_),
    .Y(_01406_)
  );
  OAI21X1 _07794_ (
    .A(execution_unit_0.inst_type_1_ ),
    .B(_01406_),
    .C(execution_unit_0.alu_0.exec_cycle ),
    .Y(_01407_)
  );
  NAND2X1 _07795_ (
    .A(_01103_),
    .B(_01407_),
    .Y(execution_unit_0.reg_dest_wr )
  );
  OR2X1 _07796_ (
    .A(execution_unit_0.inst_as_1_ ),
    .B(_01299_),
    .Y(_01408_)
  );
  NOR2X1 _07797_ (
    .A(_01163_),
    .B(_01408_),
    .Y(_01409_)
  );
  NOR2X1 _07798_ (
    .A(_01301_),
    .B(_01409_),
    .Y(_01410_)
  );
  OAI21X1 _07799_ (
    .A(execution_unit_0.inst_irq_rst ),
    .B(_01113_),
    .C(_01410_),
    .Y(execution_unit_0.reg_sp_wr )
  );
  OAI21X1 _07800_ (
    .A(_01070_),
    .B(_01106_),
    .C(_01286_),
    .Y(execution_unit_0.reg_pc_call )
  );
  AOI22X1 _07801_ (
    .A(execution_unit_0.inst_as_3_ ),
    .B(exec_done),
    .C(execution_unit_0.alu_0.exec_cycle ),
    .D(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .Y(_01411_)
  );
  OAI21X1 _07802_ (
    .A(_01066_),
    .B(_01110_),
    .C(_01411_),
    .Y(execution_unit_0.reg_incr )
  );
  AOI21X1 _07803_ (
    .A(dbg_0.UNUSED_eu_mab_0_ ),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01119_),
    .Y(dbg_0.UNUSED_eu_mb_wr_0_ )
  );
  AOI21X1 _07804_ (
    .A(_01069_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01119_),
    .Y(dbg_0.UNUSED_eu_mb_wr_1_ )
  );
  DFFSR _07805_ (
    .CLK(dco_clk),
    .D(_01029_),
    .Q(execution_unit_0.mdb_in_buf_0_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07806_ (
    .CLK(dco_clk),
    .D(_01036_),
    .Q(execution_unit_0.mdb_in_buf_1_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07807_ (
    .CLK(dco_clk),
    .D(_01037_),
    .Q(execution_unit_0.mdb_in_buf_2_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07808_ (
    .CLK(dco_clk),
    .D(_01038_),
    .Q(execution_unit_0.mdb_in_buf_3_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07809_ (
    .CLK(dco_clk),
    .D(_01039_),
    .Q(execution_unit_0.mdb_in_buf_4_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07810_ (
    .CLK(dco_clk),
    .D(_01040_),
    .Q(execution_unit_0.mdb_in_buf_5_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07811_ (
    .CLK(dco_clk),
    .D(_01041_),
    .Q(execution_unit_0.mdb_in_buf_6_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07812_ (
    .CLK(dco_clk),
    .D(_01042_),
    .Q(execution_unit_0.mdb_in_buf_7_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07813_ (
    .CLK(dco_clk),
    .D(_01043_),
    .Q(execution_unit_0.mdb_in_buf_8_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07814_ (
    .CLK(dco_clk),
    .D(_01044_),
    .Q(execution_unit_0.mdb_in_buf_9_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07815_ (
    .CLK(dco_clk),
    .D(_01030_),
    .Q(execution_unit_0.mdb_in_buf_10_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07816_ (
    .CLK(dco_clk),
    .D(_01031_),
    .Q(execution_unit_0.mdb_in_buf_11_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07817_ (
    .CLK(dco_clk),
    .D(_01032_),
    .Q(execution_unit_0.mdb_in_buf_12_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07818_ (
    .CLK(dco_clk),
    .D(_01033_),
    .Q(execution_unit_0.mdb_in_buf_13_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07819_ (
    .CLK(dco_clk),
    .D(_01034_),
    .Q(execution_unit_0.mdb_in_buf_14_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07820_ (
    .CLK(dco_clk),
    .D(_01035_),
    .Q(execution_unit_0.mdb_in_buf_15_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07821_ (
    .CLK(dco_clk),
    .D(_01046_),
    .Q(execution_unit_0.mdb_in_buf_valid ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07822_ (
    .CLK(dco_clk),
    .D(_01045_),
    .Q(execution_unit_0.mdb_in_buf_en ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07823_ (
    .CLK(dco_clk),
    .D(_01028_),
    .Q(execution_unit_0.mab_lsb ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07824_ (
    .CLK(dco_clk),
    .D(_01047_),
    .Q(eu_mdb_out_0_),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07825_ (
    .CLK(dco_clk),
    .D(_01054_),
    .Q(eu_mdb_out_1_),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07826_ (
    .CLK(dco_clk),
    .D(_01055_),
    .Q(eu_mdb_out_2_),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07827_ (
    .CLK(dco_clk),
    .D(_01056_),
    .Q(eu_mdb_out_3_),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07828_ (
    .CLK(dco_clk),
    .D(_01057_),
    .Q(eu_mdb_out_4_),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07829_ (
    .CLK(dco_clk),
    .D(_01058_),
    .Q(eu_mdb_out_5_),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07830_ (
    .CLK(dco_clk),
    .D(_01059_),
    .Q(eu_mdb_out_6_),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07831_ (
    .CLK(dco_clk),
    .D(_01060_),
    .Q(eu_mdb_out_7_),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07832_ (
    .CLK(dco_clk),
    .D(_01061_),
    .Q(execution_unit_0.mdb_out_nxt_8_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07833_ (
    .CLK(dco_clk),
    .D(_01062_),
    .Q(execution_unit_0.mdb_out_nxt_9_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07834_ (
    .CLK(dco_clk),
    .D(_01048_),
    .Q(execution_unit_0.mdb_out_nxt_10_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07835_ (
    .CLK(dco_clk),
    .D(_01049_),
    .Q(execution_unit_0.mdb_out_nxt_11_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07836_ (
    .CLK(dco_clk),
    .D(_01050_),
    .Q(execution_unit_0.mdb_out_nxt_12_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07837_ (
    .CLK(dco_clk),
    .D(_01051_),
    .Q(execution_unit_0.mdb_out_nxt_13_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07838_ (
    .CLK(dco_clk),
    .D(_01052_),
    .Q(execution_unit_0.mdb_out_nxt_14_ ),
    .R(_01063_),
    .S(1'h1)
  );
  DFFSR _07839_ (
    .CLK(dco_clk),
    .D(_01053_),
    .Q(execution_unit_0.mdb_out_nxt_15_ ),
    .R(_01063_),
    .S(1'h1)
  );
  INVX1 _07840_ (
    .A(execution_unit_0.alu_0.exec_cycle ),
    .Y(_01957_)
  );
  INVX1 _07841_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .Y(_01412_)
  );
  INVX1 _07842_ (
    .A(execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01413_)
  );
  INVX1 _07843_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_01414_)
  );
  INVX1 _07844_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01415_)
  );
  INVX1 _07845_ (
    .A(execution_unit_0.alu_0.status_0_ ),
    .Y(_01416_)
  );
  INVX1 _07846_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01417_)
  );
  INVX1 _07847_ (
    .A(execution_unit_0.alu_0.inst_jmp_4_ ),
    .Y(_01418_)
  );
  INVX1 _07848_ (
    .A(execution_unit_0.alu_0.inst_jmp_1_ ),
    .Y(_01419_)
  );
  INVX1 _07849_ (
    .A(execution_unit_0.alu_0.alu_shift_3_ ),
    .Y(_01420_)
  );
  INVX1 _07850_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .Y(_01421_)
  );
  INVX1 _07851_ (
    .A(execution_unit_0.alu_0.op_dst_15_ ),
    .Y(_01422_)
  );
  OR2X1 _07852_ (
    .A(cpu_halt_st),
    .B(execution_unit_0.alu_0.inst_so_7_ ),
    .Y(_01423_)
  );
  NOR2X1 _07853_ (
    .A(execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01423_),
    .Y(_01424_)
  );
  OR2X1 _07854_ (
    .A(execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01423_),
    .Y(_01425_)
  );
  AND2X1 _07855_ (
    .A(execution_unit_0.alu_0.inst_alu_0_ ),
    .B(execution_unit_0.alu_0.exec_cycle ),
    .Y(_01426_)
  );
  NAND2X1 _07856_ (
    .A(execution_unit_0.alu_0.inst_alu_0_ ),
    .B(execution_unit_0.alu_0.exec_cycle ),
    .Y(_01427_)
  );
  XNOR2X1 _07857_ (
    .A(execution_unit_0.alu_0.alu_swpb_8_ ),
    .B(_01427_),
    .Y(_01428_)
  );
  AND2X1 _07858_ (
    .A(execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01428_),
    .Y(_01429_)
  );
  NAND2X1 _07859_ (
    .A(execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01428_),
    .Y(_01430_)
  );
  NAND2X1 _07860_ (
    .A(execution_unit_0.alu_0.status_1_ ),
    .B(execution_unit_0.alu_0.inst_jmp_0_ ),
    .Y(_01431_)
  );
  OAI21X1 _07861_ (
    .A(_01419_),
    .B(execution_unit_0.alu_0.status_1_ ),
    .C(_01431_),
    .Y(_01432_)
  );
  MUX2X1 _07862_ (
    .A(execution_unit_0.alu_0.inst_jmp_2_ ),
    .B(execution_unit_0.alu_0.inst_jmp_3_ ),
    .S(execution_unit_0.alu_0.status_0_ ),
    .Y(_01433_)
  );
  OAI21X1 _07863_ (
    .A(execution_unit_0.alu_0.status_2_ ),
    .B(_01418_),
    .C(_01433_),
    .Y(_01434_)
  );
  NOR2X1 _07864_ (
    .A(_01432_),
    .B(_01434_),
    .Y(_01435_)
  );
  XOR2X1 _07865_ (
    .A(execution_unit_0.alu_0.status_3_ ),
    .B(execution_unit_0.alu_0.status_2_ ),
    .Y(_01436_)
  );
  MUX2X1 _07866_ (
    .A(execution_unit_0.alu_0.inst_jmp_5_ ),
    .B(execution_unit_0.alu_0.inst_jmp_6_ ),
    .S(_01436_),
    .Y(_01437_)
  );
  AND2X1 _07867_ (
    .A(_01435_),
    .B(_01437_),
    .Y(_01438_)
  );
  NAND2X1 _07868_ (
    .A(_01435_),
    .B(_01437_),
    .Y(_01439_)
  );
  AOI21X1 _07869_ (
    .A(_01428_),
    .B(_01438_),
    .C(execution_unit_0.alu_0.op_dst_0_ ),
    .Y(_01440_)
  );
  AOI21X1 _07870_ (
    .A(_01429_),
    .B(_01438_),
    .C(_01440_),
    .Y(dbg_0.UNUSED_eu_mab_0_ )
  );
  AOI21X1 _07871_ (
    .A(execution_unit_0.alu_0.status_0_ ),
    .B(execution_unit_0.alu_0.inst_alu_2_ ),
    .C(execution_unit_0.alu_0.inst_alu_1_ ),
    .Y(_01441_)
  );
  NOR2X1 _07872_ (
    .A(_01957_),
    .B(_01441_),
    .Y(_01442_)
  );
  NAND2X1 _07873_ (
    .A(dbg_0.UNUSED_eu_mab_0_ ),
    .B(_01442_),
    .Y(_01443_)
  );
  OR2X1 _07874_ (
    .A(dbg_0.UNUSED_eu_mab_0_ ),
    .B(_01442_),
    .Y(_01444_)
  );
  NOR2X1 _07875_ (
    .A(execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01428_),
    .Y(_01445_)
  );
  OR2X1 _07876_ (
    .A(execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01428_),
    .Y(_01446_)
  );
  NAND2X1 _07877_ (
    .A(_01430_),
    .B(_01446_),
    .Y(_01447_)
  );
  XNOR2X1 _07878_ (
    .A(execution_unit_0.alu_0.status_0_ ),
    .B(_01447_),
    .Y(_01448_)
  );
  NOR2X1 _07879_ (
    .A(execution_unit_0.alu_0.inst_alu_5_ ),
    .B(execution_unit_0.alu_0.inst_so_3_ ),
    .Y(_01449_)
  );
  NOR2X1 _07880_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_01450_)
  );
  NAND2X1 _07881_ (
    .A(_01415_),
    .B(_01450_),
    .Y(_01451_)
  );
  NAND2X1 _07882_ (
    .A(_01412_),
    .B(_01449_),
    .Y(_01452_)
  );
  NOR2X1 _07883_ (
    .A(_01451_),
    .B(_01452_),
    .Y(_01453_)
  );
  AOI21X1 _07884_ (
    .A(execution_unit_0.alu_0.alu_shift_0_ ),
    .B(execution_unit_0.alu_0.inst_alu_10_ ),
    .C(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01454_)
  );
  AOI22X1 _07885_ (
    .A(execution_unit_0.alu_0.alu_swpb_0_ ),
    .B(execution_unit_0.alu_0.inst_so_1_ ),
    .C(execution_unit_0.alu_0.inst_so_3_ ),
    .D(execution_unit_0.alu_0.alu_swpb_8_ ),
    .Y(_01455_)
  );
  NAND2X1 _07886_ (
    .A(_01454_),
    .B(_01455_),
    .Y(_01456_)
  );
  AOI21X1 _07887_ (
    .A(_01428_),
    .B(_01453_),
    .C(_01456_),
    .Y(_01457_)
  );
  OAI21X1 _07888_ (
    .A(_01414_),
    .B(_01430_),
    .C(_01457_),
    .Y(_01458_)
  );
  AOI21X1 _07889_ (
    .A(execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_01446_),
    .C(_01458_),
    .Y(_01459_)
  );
  OAI21X1 _07890_ (
    .A(_01412_),
    .B(_01447_),
    .C(_01459_),
    .Y(_01460_)
  );
  OAI21X1 _07891_ (
    .A(_01417_),
    .B(_01448_),
    .C(_01460_),
    .Y(_01461_)
  );
  NAND3X1 _07892_ (
    .A(_01425_),
    .B(_01443_),
    .C(_01444_),
    .Y(_01462_)
  );
  OAI21X1 _07893_ (
    .A(_01425_),
    .B(_01461_),
    .C(_01462_),
    .Y(execution_unit_0.alu_0.alu_out_0_ )
  );
  XNOR2X1 _07894_ (
    .A(execution_unit_0.alu_0.alu_shift_0_ ),
    .B(_01427_),
    .Y(_01463_)
  );
  AND2X1 _07895_ (
    .A(execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01463_),
    .Y(_01464_)
  );
  NAND2X1 _07896_ (
    .A(execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01463_),
    .Y(_01465_)
  );
  NOR2X1 _07897_ (
    .A(execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01463_),
    .Y(_01466_)
  );
  NOR2X1 _07898_ (
    .A(_01464_),
    .B(_01466_),
    .Y(_01467_)
  );
  OR2X1 _07899_ (
    .A(_01464_),
    .B(_01466_),
    .Y(_01468_)
  );
  NAND3X1 _07900_ (
    .A(_01429_),
    .B(_01438_),
    .C(_01467_),
    .Y(_01469_)
  );
  NAND3X1 _07901_ (
    .A(_01430_),
    .B(_01438_),
    .C(_01468_),
    .Y(_01470_)
  );
  AND2X1 _07902_ (
    .A(_01469_),
    .B(_01470_),
    .Y(_01471_)
  );
  OAI21X1 _07903_ (
    .A(execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01438_),
    .C(_01471_),
    .Y(_01472_)
  );
  INVX1 _07904_ (
    .A(_01472_),
    .Y(dbg_0.UNUSED_eu_mab_1_ )
  );
  OR2X1 _07905_ (
    .A(_01443_),
    .B(_01472_),
    .Y(_01473_)
  );
  OAI21X1 _07906_ (
    .A(_01443_),
    .B(_01472_),
    .C(_01425_),
    .Y(_01474_)
  );
  AOI21X1 _07907_ (
    .A(_01443_),
    .B(_01472_),
    .C(_01474_),
    .Y(_01475_)
  );
  AOI21X1 _07908_ (
    .A(execution_unit_0.alu_0.status_0_ ),
    .B(_01446_),
    .C(_01429_),
    .Y(_01476_)
  );
  OAI21X1 _07909_ (
    .A(_01416_),
    .B(_01445_),
    .C(_01430_),
    .Y(_01477_)
  );
  XNOR2X1 _07910_ (
    .A(_01468_),
    .B(_01476_),
    .Y(_01478_)
  );
  INVX1 _07911_ (
    .A(_01478_),
    .Y(_01479_)
  );
  AOI21X1 _07912_ (
    .A(_01467_),
    .B(_01477_),
    .C(_01464_),
    .Y(_01480_)
  );
  OAI21X1 _07913_ (
    .A(_01468_),
    .B(_01476_),
    .C(_01465_),
    .Y(_01481_)
  );
  XNOR2X1 _07914_ (
    .A(execution_unit_0.alu_0.alu_shift_1_ ),
    .B(_01427_),
    .Y(_01482_)
  );
  AND2X1 _07915_ (
    .A(execution_unit_0.alu_0.op_dst_2_ ),
    .B(_01482_),
    .Y(_01483_)
  );
  NAND2X1 _07916_ (
    .A(execution_unit_0.alu_0.op_dst_2_ ),
    .B(_01482_),
    .Y(_01484_)
  );
  OR2X1 _07917_ (
    .A(execution_unit_0.alu_0.op_dst_2_ ),
    .B(_01482_),
    .Y(_01485_)
  );
  INVX1 _07918_ (
    .A(_01485_),
    .Y(_01486_)
  );
  NAND2X1 _07919_ (
    .A(_01484_),
    .B(_01485_),
    .Y(_01487_)
  );
  XNOR2X1 _07920_ (
    .A(_01481_),
    .B(_01487_),
    .Y(_01488_)
  );
  NOR2X1 _07921_ (
    .A(_01479_),
    .B(_01488_),
    .Y(_01489_)
  );
  OR2X1 _07922_ (
    .A(_01479_),
    .B(_01488_),
    .Y(_01490_)
  );
  AOI21X1 _07923_ (
    .A(_01481_),
    .B(_01485_),
    .C(_01483_),
    .Y(_01491_)
  );
  OAI21X1 _07924_ (
    .A(_01480_),
    .B(_01486_),
    .C(_01484_),
    .Y(_01492_)
  );
  XNOR2X1 _07925_ (
    .A(execution_unit_0.alu_0.alu_shift_2_ ),
    .B(_01427_),
    .Y(_01493_)
  );
  AND2X1 _07926_ (
    .A(execution_unit_0.alu_0.op_dst_3_ ),
    .B(_01493_),
    .Y(_01494_)
  );
  NAND2X1 _07927_ (
    .A(execution_unit_0.alu_0.op_dst_3_ ),
    .B(_01493_),
    .Y(_01495_)
  );
  OR2X1 _07928_ (
    .A(execution_unit_0.alu_0.op_dst_3_ ),
    .B(_01493_),
    .Y(_01496_)
  );
  INVX1 _07929_ (
    .A(_01496_),
    .Y(_01497_)
  );
  NAND2X1 _07930_ (
    .A(_01495_),
    .B(_01496_),
    .Y(_01498_)
  );
  XNOR2X1 _07931_ (
    .A(_01492_),
    .B(_01498_),
    .Y(_01499_)
  );
  XNOR2X1 _07932_ (
    .A(_01491_),
    .B(_01498_),
    .Y(_01500_)
  );
  OAI21X1 _07933_ (
    .A(_01492_),
    .B(_01494_),
    .C(_01496_),
    .Y(_01501_)
  );
  AOI21X1 _07934_ (
    .A(_01491_),
    .B(_01495_),
    .C(_01497_),
    .Y(_01502_)
  );
  AOI21X1 _07935_ (
    .A(_01490_),
    .B(_01499_),
    .C(_01502_),
    .Y(_01503_)
  );
  OAI21X1 _07936_ (
    .A(_01489_),
    .B(_01500_),
    .C(_01501_),
    .Y(_01504_)
  );
  NAND2X1 _07937_ (
    .A(_01478_),
    .B(_01504_),
    .Y(_01505_)
  );
  AOI21X1 _07938_ (
    .A(_01479_),
    .B(_01503_),
    .C(_01417_),
    .Y(_01506_)
  );
  OAI21X1 _07939_ (
    .A(execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01463_),
    .C(execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01507_)
  );
  NAND2X1 _07940_ (
    .A(_01453_),
    .B(_01463_),
    .Y(_01508_)
  );
  AOI22X1 _07941_ (
    .A(execution_unit_0.alu_0.alu_shift_0_ ),
    .B(execution_unit_0.alu_0.inst_so_3_ ),
    .C(_01464_),
    .D(execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_01509_)
  );
  OAI21X1 _07942_ (
    .A(_01412_),
    .B(_01468_),
    .C(_01509_),
    .Y(_01510_)
  );
  AOI22X1 _07943_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_8_ ),
    .C(execution_unit_0.alu_0.alu_shift_1_ ),
    .D(execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01511_)
  );
  NAND3X1 _07944_ (
    .A(_01507_),
    .B(_01508_),
    .C(_01511_),
    .Y(_01512_)
  );
  OR2X1 _07945_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01512_),
    .Y(_01513_)
  );
  OAI21X1 _07946_ (
    .A(_01510_),
    .B(_01513_),
    .C(_01424_),
    .Y(_01514_)
  );
  AOI21X1 _07947_ (
    .A(_01505_),
    .B(_01506_),
    .C(_01514_),
    .Y(_01515_)
  );
  NOR2X1 _07948_ (
    .A(_01475_),
    .B(_01515_),
    .Y(_01516_)
  );
  INVX1 _07949_ (
    .A(_01516_),
    .Y(execution_unit_0.alu_0.alu_out_1_ )
  );
  OAI21X1 _07950_ (
    .A(_01439_),
    .B(_01465_),
    .C(_01469_),
    .Y(_01517_)
  );
  AOI21X1 _07951_ (
    .A(_01438_),
    .B(_01482_),
    .C(execution_unit_0.alu_0.op_dst_2_ ),
    .Y(_01518_)
  );
  AOI21X1 _07952_ (
    .A(_01438_),
    .B(_01483_),
    .C(_01518_),
    .Y(_01519_)
  );
  XNOR2X1 _07953_ (
    .A(_01517_),
    .B(_01519_),
    .Y(_01520_)
  );
  INVX1 _07954_ (
    .A(_01520_),
    .Y(dbg_0.UNUSED_eu_mab_2_ )
  );
  AND2X1 _07955_ (
    .A(_01473_),
    .B(_01520_),
    .Y(_01521_)
  );
  NOR2X1 _07956_ (
    .A(_01473_),
    .B(_01520_),
    .Y(_01522_)
  );
  OAI21X1 _07957_ (
    .A(_01473_),
    .B(_01520_),
    .C(_01425_),
    .Y(_01523_)
  );
  OAI21X1 _07958_ (
    .A(_01490_),
    .B(_01501_),
    .C(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01524_)
  );
  AOI21X1 _07959_ (
    .A(_01488_),
    .B(_01505_),
    .C(_01524_),
    .Y(_01525_)
  );
  AOI22X1 _07960_ (
    .A(execution_unit_0.alu_0.inst_so_3_ ),
    .B(execution_unit_0.alu_0.alu_shift_1_ ),
    .C(execution_unit_0.alu_0.alu_shift_2_ ),
    .D(execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01526_)
  );
  OAI21X1 _07961_ (
    .A(_01414_),
    .B(_01484_),
    .C(_01526_),
    .Y(_01527_)
  );
  AOI21X1 _07962_ (
    .A(_01453_),
    .B(_01482_),
    .C(execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01528_)
  );
  NOR2X1 _07963_ (
    .A(_01486_),
    .B(_01528_),
    .Y(_01529_)
  );
  OR2X1 _07964_ (
    .A(_01527_),
    .B(_01529_),
    .Y(_01530_)
  );
  AOI21X1 _07965_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_9_ ),
    .C(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01531_)
  );
  OAI21X1 _07966_ (
    .A(_01412_),
    .B(_01487_),
    .C(_01531_),
    .Y(_01532_)
  );
  OAI21X1 _07967_ (
    .A(_01530_),
    .B(_01532_),
    .C(_01424_),
    .Y(_01533_)
  );
  OAI22X1 _07968_ (
    .A(_01521_),
    .B(_01523_),
    .C(_01525_),
    .D(_01533_),
    .Y(execution_unit_0.alu_0.alu_out_2_ )
  );
  AOI22X1 _07969_ (
    .A(_01438_),
    .B(_01483_),
    .C(_01517_),
    .D(_01519_),
    .Y(_01534_)
  );
  OAI21X1 _07970_ (
    .A(execution_unit_0.alu_0.op_dst_3_ ),
    .B(_01438_),
    .C(_01496_),
    .Y(_01535_)
  );
  AOI21X1 _07971_ (
    .A(_01438_),
    .B(_01494_),
    .C(_01535_),
    .Y(_01536_)
  );
  XNOR2X1 _07972_ (
    .A(_01534_),
    .B(_01536_),
    .Y(dbg_0.UNUSED_eu_mab_3_ )
  );
  NAND2X1 _07973_ (
    .A(_01522_),
    .B(dbg_0.UNUSED_eu_mab_3_ ),
    .Y(_01537_)
  );
  XNOR2X1 _07974_ (
    .A(_01522_),
    .B(dbg_0.UNUSED_eu_mab_3_ ),
    .Y(_01538_)
  );
  OAI21X1 _07975_ (
    .A(_01489_),
    .B(_01501_),
    .C(_01500_),
    .Y(_01539_)
  );
  AND2X1 _07976_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01539_),
    .Y(_01540_)
  );
  OAI21X1 _07977_ (
    .A(_01489_),
    .B(_01500_),
    .C(_01540_),
    .Y(_01541_)
  );
  NAND2X1 _07978_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01424_),
    .Y(_01542_)
  );
  AOI22X1 _07979_ (
    .A(execution_unit_0.alu_0.inst_so_3_ ),
    .B(execution_unit_0.alu_0.alu_shift_2_ ),
    .C(execution_unit_0.alu_0.alu_shift_10_ ),
    .D(execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01543_)
  );
  OAI21X1 _07980_ (
    .A(_01415_),
    .B(_01420_),
    .C(_01543_),
    .Y(_01544_)
  );
  AOI22X1 _07981_ (
    .A(_01453_),
    .B(_01493_),
    .C(_01496_),
    .D(execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01545_)
  );
  AOI21X1 _07982_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01494_),
    .C(_01544_),
    .Y(_01546_)
  );
  NAND2X1 _07983_ (
    .A(_01545_),
    .B(_01546_),
    .Y(_01547_)
  );
  OAI21X1 _07984_ (
    .A(_01412_),
    .B(_01498_),
    .C(_01424_),
    .Y(_01548_)
  );
  OAI21X1 _07985_ (
    .A(_01547_),
    .B(_01548_),
    .C(_01542_),
    .Y(_01549_)
  );
  AOI22X1 _07986_ (
    .A(_01425_),
    .B(_01538_),
    .C(_01541_),
    .D(_01549_),
    .Y(execution_unit_0.alu_0.alu_out_3_ )
  );
  XNOR2X1 _07987_ (
    .A(_01420_),
    .B(_01426_),
    .Y(_01550_)
  );
  AND2X1 _07988_ (
    .A(execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01550_),
    .Y(_01551_)
  );
  NAND2X1 _07989_ (
    .A(execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01550_),
    .Y(_01552_)
  );
  NAND2X1 _07990_ (
    .A(_01438_),
    .B(_01550_),
    .Y(_01553_)
  );
  XOR2X1 _07991_ (
    .A(execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01553_),
    .Y(_01554_)
  );
  INVX1 _07992_ (
    .A(_01554_),
    .Y(_01555_)
  );
  OAI22X1 _07993_ (
    .A(_01439_),
    .B(_01495_),
    .C(_01534_),
    .D(_01535_),
    .Y(_01556_)
  );
  XNOR2X1 _07994_ (
    .A(_01555_),
    .B(_01556_),
    .Y(_01557_)
  );
  INVX1 _07995_ (
    .A(_01557_),
    .Y(dbg_0.UNUSED_eu_mab_4_ )
  );
  AND2X1 _07996_ (
    .A(_01537_),
    .B(_01557_),
    .Y(_01558_)
  );
  NOR2X1 _07997_ (
    .A(_01537_),
    .B(_01557_),
    .Y(_01559_)
  );
  NOR2X1 _07998_ (
    .A(execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01550_),
    .Y(_01560_)
  );
  NOR2X1 _07999_ (
    .A(_01551_),
    .B(_01560_),
    .Y(_01561_)
  );
  OR2X1 _08000_ (
    .A(_01551_),
    .B(_01560_),
    .Y(_01562_)
  );
  NOR3X1 _08001_ (
    .A(_01489_),
    .B(_01500_),
    .C(_01501_),
    .Y(_01563_)
  );
  NAND3X1 _08002_ (
    .A(_01490_),
    .B(_01499_),
    .C(_01502_),
    .Y(_01564_)
  );
  NOR3X1 _08003_ (
    .A(_01503_),
    .B(_01562_),
    .C(_01563_),
    .Y(_01565_)
  );
  NAND3X1 _08004_ (
    .A(_01504_),
    .B(_01561_),
    .C(_01564_),
    .Y(_01566_)
  );
  AOI21X1 _08005_ (
    .A(_01504_),
    .B(_01564_),
    .C(_01561_),
    .Y(_01567_)
  );
  OAI21X1 _08006_ (
    .A(_01565_),
    .B(_01567_),
    .C(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01568_)
  );
  NOR2X1 _08007_ (
    .A(_01413_),
    .B(_01560_),
    .Y(_01569_)
  );
  AOI21X1 _08008_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_4_ ),
    .C(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01570_)
  );
  AOI22X1 _08009_ (
    .A(execution_unit_0.alu_0.inst_so_3_ ),
    .B(execution_unit_0.alu_0.alu_shift_3_ ),
    .C(execution_unit_0.alu_0.alu_shift_11_ ),
    .D(execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01571_)
  );
  NAND2X1 _08010_ (
    .A(_01570_),
    .B(_01571_),
    .Y(_01572_)
  );
  AOI21X1 _08011_ (
    .A(_01453_),
    .B(_01550_),
    .C(_01572_),
    .Y(_01573_)
  );
  OAI21X1 _08012_ (
    .A(_01414_),
    .B(_01552_),
    .C(_01573_),
    .Y(_01574_)
  );
  NOR2X1 _08013_ (
    .A(_01569_),
    .B(_01574_),
    .Y(_01575_)
  );
  OAI21X1 _08014_ (
    .A(_01412_),
    .B(_01562_),
    .C(_01575_),
    .Y(_01576_)
  );
  OAI21X1 _08015_ (
    .A(_01537_),
    .B(_01557_),
    .C(_01425_),
    .Y(_01577_)
  );
  NAND3X1 _08016_ (
    .A(_01424_),
    .B(_01568_),
    .C(_01576_),
    .Y(_01578_)
  );
  OAI21X1 _08017_ (
    .A(_01558_),
    .B(_01577_),
    .C(_01578_),
    .Y(execution_unit_0.alu_0.alu_out_4_ )
  );
  AOI22X1 _08018_ (
    .A(_01438_),
    .B(_01551_),
    .C(_01555_),
    .D(_01556_),
    .Y(_01579_)
  );
  XNOR2X1 _08019_ (
    .A(execution_unit_0.alu_0.alu_shift_4_ ),
    .B(_01427_),
    .Y(_01580_)
  );
  AND2X1 _08020_ (
    .A(execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01580_),
    .Y(_01581_)
  );
  NAND2X1 _08021_ (
    .A(execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01580_),
    .Y(_01582_)
  );
  NAND2X1 _08022_ (
    .A(_01438_),
    .B(_01580_),
    .Y(_01583_)
  );
  XOR2X1 _08023_ (
    .A(execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01583_),
    .Y(_01584_)
  );
  XOR2X1 _08024_ (
    .A(_01579_),
    .B(_01584_),
    .Y(dbg_0.UNUSED_eu_mab_5_ )
  );
  NOR2X1 _08025_ (
    .A(_01559_),
    .B(dbg_0.UNUSED_eu_mab_5_ ),
    .Y(_01585_)
  );
  NAND2X1 _08026_ (
    .A(_01559_),
    .B(dbg_0.UNUSED_eu_mab_5_ ),
    .Y(_01586_)
  );
  OAI21X1 _08027_ (
    .A(execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01423_),
    .C(_01586_),
    .Y(_01587_)
  );
  XNOR2X1 _08028_ (
    .A(execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01580_),
    .Y(_01588_)
  );
  INVX1 _08029_ (
    .A(_01588_),
    .Y(_01589_)
  );
  AOI21X1 _08030_ (
    .A(_01552_),
    .B(_01566_),
    .C(_01588_),
    .Y(_01590_)
  );
  OAI21X1 _08031_ (
    .A(_01551_),
    .B(_01565_),
    .C(_01589_),
    .Y(_01591_)
  );
  NAND3X1 _08032_ (
    .A(_01552_),
    .B(_01566_),
    .C(_01588_),
    .Y(_01592_)
  );
  AND2X1 _08033_ (
    .A(_01591_),
    .B(_01592_),
    .Y(_01593_)
  );
  XNOR2X1 _08034_ (
    .A(execution_unit_0.alu_0.alu_shift_5_ ),
    .B(_01427_),
    .Y(_01594_)
  );
  AND2X1 _08035_ (
    .A(execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01594_),
    .Y(_01595_)
  );
  NAND2X1 _08036_ (
    .A(execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01594_),
    .Y(_01596_)
  );
  XNOR2X1 _08037_ (
    .A(execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01594_),
    .Y(_01597_)
  );
  INVX1 _08038_ (
    .A(_01597_),
    .Y(_01598_)
  );
  AOI21X1 _08039_ (
    .A(_01582_),
    .B(_01591_),
    .C(_01597_),
    .Y(_01599_)
  );
  OAI21X1 _08040_ (
    .A(_01581_),
    .B(_01590_),
    .C(_01598_),
    .Y(_01600_)
  );
  NAND3X1 _08041_ (
    .A(_01582_),
    .B(_01591_),
    .C(_01597_),
    .Y(_01601_)
  );
  NAND2X1 _08042_ (
    .A(_01600_),
    .B(_01601_),
    .Y(_01602_)
  );
  AOI21X1 _08043_ (
    .A(_01600_),
    .B(_01601_),
    .C(_01593_),
    .Y(_01603_)
  );
  XNOR2X1 _08044_ (
    .A(execution_unit_0.alu_0.alu_shift_6_ ),
    .B(_01427_),
    .Y(_01604_)
  );
  AND2X1 _08045_ (
    .A(execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01604_),
    .Y(_01605_)
  );
  NOR2X1 _08046_ (
    .A(execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01604_),
    .Y(_01606_)
  );
  NOR2X1 _08047_ (
    .A(_01605_),
    .B(_01606_),
    .Y(_01607_)
  );
  INVX1 _08048_ (
    .A(_01607_),
    .Y(_01608_)
  );
  NAND3X1 _08049_ (
    .A(_01596_),
    .B(_01600_),
    .C(_01607_),
    .Y(_01609_)
  );
  OAI21X1 _08050_ (
    .A(_01595_),
    .B(_01599_),
    .C(_01608_),
    .Y(_01610_)
  );
  NAND2X1 _08051_ (
    .A(_01609_),
    .B(_01610_),
    .Y(_01611_)
  );
  AOI21X1 _08052_ (
    .A(_01609_),
    .B(_01610_),
    .C(_01603_),
    .Y(_01612_)
  );
  INVX1 _08053_ (
    .A(_01612_),
    .Y(_01613_)
  );
  AOI21X1 _08054_ (
    .A(_01596_),
    .B(_01600_),
    .C(_01606_),
    .Y(_01614_)
  );
  NOR2X1 _08055_ (
    .A(_01605_),
    .B(_01614_),
    .Y(_01615_)
  );
  NAND2X1 _08056_ (
    .A(_01613_),
    .B(_01615_),
    .Y(_01616_)
  );
  AOI21X1 _08057_ (
    .A(_01613_),
    .B(_01615_),
    .C(_01593_),
    .Y(_01617_)
  );
  XNOR2X1 _08058_ (
    .A(_01593_),
    .B(_01616_),
    .Y(_01618_)
  );
  NOR2X1 _08059_ (
    .A(_01412_),
    .B(_01588_),
    .Y(_01619_)
  );
  OAI21X1 _08060_ (
    .A(execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01580_),
    .C(execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01620_)
  );
  NAND2X1 _08061_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01581_),
    .Y(_01621_)
  );
  AOI21X1 _08062_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_5_ ),
    .C(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01622_)
  );
  AOI22X1 _08063_ (
    .A(execution_unit_0.alu_0.inst_so_3_ ),
    .B(execution_unit_0.alu_0.alu_shift_4_ ),
    .C(execution_unit_0.alu_0.alu_shift_12_ ),
    .D(execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01623_)
  );
  NAND2X1 _08064_ (
    .A(_01622_),
    .B(_01623_),
    .Y(_01624_)
  );
  AOI21X1 _08065_ (
    .A(_01453_),
    .B(_01580_),
    .C(_01624_),
    .Y(_01625_)
  );
  NAND3X1 _08066_ (
    .A(_01620_),
    .B(_01621_),
    .C(_01625_),
    .Y(_01626_)
  );
  OAI21X1 _08067_ (
    .A(_01619_),
    .B(_01626_),
    .C(_01424_),
    .Y(_01627_)
  );
  AOI21X1 _08068_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01618_),
    .C(_01627_),
    .Y(_01628_)
  );
  INVX1 _08069_ (
    .A(_01628_),
    .Y(_01629_)
  );
  OAI21X1 _08070_ (
    .A(_01585_),
    .B(_01587_),
    .C(_01629_),
    .Y(execution_unit_0.alu_0.alu_out_5_ )
  );
  OAI22X1 _08071_ (
    .A(_01439_),
    .B(_01582_),
    .C(_01584_),
    .D(_01579_),
    .Y(_01630_)
  );
  NAND2X1 _08072_ (
    .A(_01438_),
    .B(_01594_),
    .Y(_01631_)
  );
  XOR2X1 _08073_ (
    .A(execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01631_),
    .Y(_01632_)
  );
  INVX1 _08074_ (
    .A(_01632_),
    .Y(_01633_)
  );
  NAND2X1 _08075_ (
    .A(_01630_),
    .B(_01633_),
    .Y(_01634_)
  );
  XNOR2X1 _08076_ (
    .A(_01630_),
    .B(_01633_),
    .Y(_01635_)
  );
  INVX1 _08077_ (
    .A(_01635_),
    .Y(dbg_0.UNUSED_eu_mab_6_ )
  );
  NOR2X1 _08078_ (
    .A(_01586_),
    .B(_01635_),
    .Y(_01636_)
  );
  XNOR2X1 _08079_ (
    .A(_01586_),
    .B(_01635_),
    .Y(_01637_)
  );
  NOR2X1 _08080_ (
    .A(_01412_),
    .B(_01597_),
    .Y(_01638_)
  );
  OAI21X1 _08081_ (
    .A(execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01594_),
    .C(execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01639_)
  );
  AOI22X1 _08082_ (
    .A(execution_unit_0.alu_0.inst_so_3_ ),
    .B(execution_unit_0.alu_0.alu_shift_5_ ),
    .C(execution_unit_0.alu_0.alu_shift_13_ ),
    .D(execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01640_)
  );
  NAND2X1 _08083_ (
    .A(_01424_),
    .B(_01640_),
    .Y(_01641_)
  );
  AOI21X1 _08084_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_6_ ),
    .C(_01641_),
    .Y(_01642_)
  );
  AOI22X1 _08085_ (
    .A(_01453_),
    .B(_01594_),
    .C(_01595_),
    .D(execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_01643_)
  );
  NAND3X1 _08086_ (
    .A(_01639_),
    .B(_01642_),
    .C(_01643_),
    .Y(_01644_)
  );
  OAI21X1 _08087_ (
    .A(_01638_),
    .B(_01644_),
    .C(_01542_),
    .Y(_01645_)
  );
  XNOR2X1 _08088_ (
    .A(_01602_),
    .B(_01617_),
    .Y(_01646_)
  );
  NAND2X1 _08089_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01646_),
    .Y(_01647_)
  );
  AOI22X1 _08090_ (
    .A(_01425_),
    .B(_01637_),
    .C(_01645_),
    .D(_01647_),
    .Y(execution_unit_0.alu_0.alu_out_6_ )
  );
  AOI21X1 _08091_ (
    .A(_01438_),
    .B(_01604_),
    .C(execution_unit_0.alu_0.op_dst_7_ ),
    .Y(_01648_)
  );
  AOI21X1 _08092_ (
    .A(_01438_),
    .B(_01605_),
    .C(_01648_),
    .Y(_01649_)
  );
  OAI21X1 _08093_ (
    .A(_01439_),
    .B(_01596_),
    .C(_01634_),
    .Y(_01650_)
  );
  XOR2X1 _08094_ (
    .A(_01649_),
    .B(_01650_),
    .Y(dbg_0.UNUSED_eu_mab_7_ )
  );
  NAND2X1 _08095_ (
    .A(_01636_),
    .B(dbg_0.UNUSED_eu_mab_7_ ),
    .Y(_01651_)
  );
  XNOR2X1 _08096_ (
    .A(_01636_),
    .B(dbg_0.UNUSED_eu_mab_7_ ),
    .Y(_01652_)
  );
  MUX2X1 _08097_ (
    .A(execution_unit_0.alu_0.alu_shift_6_ ),
    .B(execution_unit_0.alu_0.alu_shift_14_ ),
    .S(execution_unit_0.alu_0.inst_bw ),
    .Y(_01653_)
  );
  NAND2X1 _08098_ (
    .A(execution_unit_0.alu_0.status_0_ ),
    .B(execution_unit_0.alu_0.inst_so_0_ ),
    .Y(_01654_)
  );
  OAI21X1 _08099_ (
    .A(execution_unit_0.alu_0.inst_so_0_ ),
    .B(_01653_),
    .C(_01654_),
    .Y(_01655_)
  );
  NOR2X1 _08100_ (
    .A(_01421_),
    .B(_01655_),
    .Y(_01656_)
  );
  OAI21X1 _08101_ (
    .A(execution_unit_0.alu_0.alu_swpb_0_ ),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01657_)
  );
  NOR2X1 _08102_ (
    .A(_01656_),
    .B(_01657_),
    .Y(_01658_)
  );
  AND2X1 _08103_ (
    .A(execution_unit_0.alu_0.inst_so_3_ ),
    .B(execution_unit_0.alu_0.alu_shift_6_ ),
    .Y(_01659_)
  );
  AOI21X1 _08104_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_14_ ),
    .C(_01659_),
    .Y(_01660_)
  );
  AND2X1 _08105_ (
    .A(_01424_),
    .B(_01660_),
    .Y(_01661_)
  );
  AOI22X1 _08106_ (
    .A(_01453_),
    .B(_01604_),
    .C(_01605_),
    .D(execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_01662_)
  );
  OAI21X1 _08107_ (
    .A(_01413_),
    .B(_01606_),
    .C(_01661_),
    .Y(_01663_)
  );
  AOI21X1 _08108_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01607_),
    .C(_01663_),
    .Y(_01664_)
  );
  NAND2X1 _08109_ (
    .A(_01662_),
    .B(_01664_),
    .Y(_01665_)
  );
  OAI21X1 _08110_ (
    .A(_01658_),
    .B(_01665_),
    .C(_01542_),
    .Y(_01666_)
  );
  NOR2X1 _08111_ (
    .A(_01603_),
    .B(_01606_),
    .Y(_01667_)
  );
  NOR2X1 _08112_ (
    .A(_01417_),
    .B(_01612_),
    .Y(_01668_)
  );
  OAI21X1 _08113_ (
    .A(_01611_),
    .B(_01667_),
    .C(_01668_),
    .Y(_01669_)
  );
  AOI22X1 _08114_ (
    .A(_01425_),
    .B(_01652_),
    .C(_01666_),
    .D(_01669_),
    .Y(execution_unit_0.alu_0.alu_out_7_ )
  );
  OAI21X1 _08115_ (
    .A(_01595_),
    .B(_01605_),
    .C(_01438_),
    .Y(_01670_)
  );
  OAI22X1 _08116_ (
    .A(_01634_),
    .B(_01648_),
    .C(_01670_),
    .D(_01606_),
    .Y(_01671_)
  );
  NOR2X1 _08117_ (
    .A(_01957_),
    .B(_01421_),
    .Y(_01672_)
  );
  NAND2X1 _08118_ (
    .A(execution_unit_0.alu_0.exec_cycle ),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01673_)
  );
  OAI21X1 _08119_ (
    .A(execution_unit_0.alu_0.alu_swpb_0_ ),
    .B(_01426_),
    .C(_01673_),
    .Y(_01674_)
  );
  AOI21X1 _08120_ (
    .A(execution_unit_0.alu_0.alu_swpb_0_ ),
    .B(_01426_),
    .C(_01674_),
    .Y(_01675_)
  );
  AND2X1 _08121_ (
    .A(execution_unit_0.alu_0.op_dst_8_ ),
    .B(_01675_),
    .Y(_01676_)
  );
  INVX1 _08122_ (
    .A(_01676_),
    .Y(_01677_)
  );
  NAND2X1 _08123_ (
    .A(_01438_),
    .B(_01676_),
    .Y(_01678_)
  );
  AOI22X1 _08124_ (
    .A(execution_unit_0.alu_0.op_dst_8_ ),
    .B(_01673_),
    .C(_01675_),
    .D(_01438_),
    .Y(_01679_)
  );
  AOI21X1 _08125_ (
    .A(_01438_),
    .B(_01676_),
    .C(_01679_),
    .Y(_01680_)
  );
  NAND2X1 _08126_ (
    .A(_01671_),
    .B(_01680_),
    .Y(_01681_)
  );
  XNOR2X1 _08127_ (
    .A(_01671_),
    .B(_01680_),
    .Y(_01682_)
  );
  INVX1 _08128_ (
    .A(_01682_),
    .Y(dbg_0.UNUSED_eu_mab_8_ )
  );
  AOI21X1 _08129_ (
    .A(execution_unit_0.alu_0.op_dst_8_ ),
    .B(_01673_),
    .C(_01675_),
    .Y(_01683_)
  );
  NOR2X1 _08130_ (
    .A(_01676_),
    .B(_01683_),
    .Y(_01684_)
  );
  XNOR2X1 _08131_ (
    .A(_01612_),
    .B(_01615_),
    .Y(_01685_)
  );
  XOR2X1 _08132_ (
    .A(_01612_),
    .B(_01615_),
    .Y(_01686_)
  );
  XNOR2X1 _08133_ (
    .A(_01684_),
    .B(_01685_),
    .Y(_01687_)
  );
  NAND2X1 _08134_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01684_),
    .Y(_01688_)
  );
  NAND2X1 _08135_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01676_),
    .Y(_01689_)
  );
  AOI21X1 _08136_ (
    .A(execution_unit_0.alu_0.alu_swpb_8_ ),
    .B(execution_unit_0.alu_0.inst_so_1_ ),
    .C(_01659_),
    .Y(_01690_)
  );
  OAI21X1 _08137_ (
    .A(_01413_),
    .B(_01683_),
    .C(_01690_),
    .Y(_01691_)
  );
  AOI22X1 _08138_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_8_ ),
    .C(_01453_),
    .D(_01675_),
    .Y(_01692_)
  );
  NAND3X1 _08139_ (
    .A(_01688_),
    .B(_01689_),
    .C(_01692_),
    .Y(_01693_)
  );
  OAI21X1 _08140_ (
    .A(_01691_),
    .B(_01693_),
    .C(_01424_),
    .Y(_01694_)
  );
  AOI22X1 _08141_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01687_),
    .C(_01694_),
    .D(_01542_),
    .Y(_01695_)
  );
  INVX1 _08142_ (
    .A(_01695_),
    .Y(_01696_)
  );
  NOR2X1 _08143_ (
    .A(_01651_),
    .B(_01682_),
    .Y(_01697_)
  );
  XNOR2X1 _08144_ (
    .A(_01651_),
    .B(_01682_),
    .Y(_01698_)
  );
  OAI21X1 _08145_ (
    .A(_01424_),
    .B(_01698_),
    .C(_01696_),
    .Y(execution_unit_0.alu_0.alu_out_8_ )
  );
  XNOR2X1 _08146_ (
    .A(execution_unit_0.alu_0.alu_shift_8_ ),
    .B(_01426_),
    .Y(_01699_)
  );
  NOR2X1 _08147_ (
    .A(_01672_),
    .B(_01699_),
    .Y(_01700_)
  );
  AND2X1 _08148_ (
    .A(execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01700_),
    .Y(_01701_)
  );
  NAND2X1 _08149_ (
    .A(execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01700_),
    .Y(_01702_)
  );
  NOR2X1 _08150_ (
    .A(_01439_),
    .B(_01702_),
    .Y(_01703_)
  );
  AOI21X1 _08151_ (
    .A(execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01673_),
    .C(_01700_),
    .Y(_01704_)
  );
  AOI22X1 _08152_ (
    .A(execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01673_),
    .C(_01700_),
    .D(_01438_),
    .Y(_01705_)
  );
  NOR2X1 _08153_ (
    .A(_01703_),
    .B(_01705_),
    .Y(_01706_)
  );
  OAI21X1 _08154_ (
    .A(_01439_),
    .B(_01677_),
    .C(_01681_),
    .Y(_01707_)
  );
  XOR2X1 _08155_ (
    .A(_01706_),
    .B(_01707_),
    .Y(dbg_0.UNUSED_eu_mab_9_ )
  );
  NOR2X1 _08156_ (
    .A(_01697_),
    .B(dbg_0.UNUSED_eu_mab_9_ ),
    .Y(_01708_)
  );
  NAND2X1 _08157_ (
    .A(_01697_),
    .B(dbg_0.UNUSED_eu_mab_9_ ),
    .Y(_01709_)
  );
  OAI21X1 _08158_ (
    .A(execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01423_),
    .C(_01709_),
    .Y(_01710_)
  );
  NOR2X1 _08159_ (
    .A(_01701_),
    .B(_01704_),
    .Y(_01711_)
  );
  AOI21X1 _08160_ (
    .A(_01684_),
    .B(_01685_),
    .C(_01676_),
    .Y(_01712_)
  );
  OAI21X1 _08161_ (
    .A(_01683_),
    .B(_01686_),
    .C(_01677_),
    .Y(_01713_)
  );
  XNOR2X1 _08162_ (
    .A(_01711_),
    .B(_01712_),
    .Y(_01714_)
  );
  XNOR2X1 _08163_ (
    .A(execution_unit_0.alu_0.alu_shift_10_ ),
    .B(_01426_),
    .Y(_01715_)
  );
  NOR2X1 _08164_ (
    .A(_01672_),
    .B(_01715_),
    .Y(_01716_)
  );
  AND2X1 _08165_ (
    .A(execution_unit_0.alu_0.op_dst_11_ ),
    .B(_01716_),
    .Y(_01717_)
  );
  NAND2X1 _08166_ (
    .A(execution_unit_0.alu_0.op_dst_11_ ),
    .B(_01716_),
    .Y(_01718_)
  );
  AOI21X1 _08167_ (
    .A(execution_unit_0.alu_0.op_dst_11_ ),
    .B(_01673_),
    .C(_01716_),
    .Y(_01719_)
  );
  NOR2X1 _08168_ (
    .A(_01717_),
    .B(_01719_),
    .Y(_01720_)
  );
  XNOR2X1 _08169_ (
    .A(execution_unit_0.alu_0.alu_shift_9_ ),
    .B(_01426_),
    .Y(_01721_)
  );
  NOR2X1 _08170_ (
    .A(_01672_),
    .B(_01721_),
    .Y(_01722_)
  );
  OAI21X1 _08171_ (
    .A(_01957_),
    .B(_01421_),
    .C(execution_unit_0.alu_0.op_dst_10_ ),
    .Y(_01723_)
  );
  NOR2X1 _08172_ (
    .A(_01721_),
    .B(_01723_),
    .Y(_01724_)
  );
  INVX1 _08173_ (
    .A(_01724_),
    .Y(_01725_)
  );
  AOI21X1 _08174_ (
    .A(_01711_),
    .B(_01713_),
    .C(_01701_),
    .Y(_01726_)
  );
  OAI21X1 _08175_ (
    .A(_01704_),
    .B(_01712_),
    .C(_01702_),
    .Y(_01727_)
  );
  AOI21X1 _08176_ (
    .A(execution_unit_0.alu_0.op_dst_10_ ),
    .B(_01673_),
    .C(_01722_),
    .Y(_01728_)
  );
  NOR2X1 _08177_ (
    .A(_01724_),
    .B(_01728_),
    .Y(_01729_)
  );
  AOI21X1 _08178_ (
    .A(_01727_),
    .B(_01729_),
    .C(_01724_),
    .Y(_01730_)
  );
  OAI21X1 _08179_ (
    .A(_01726_),
    .B(_01728_),
    .C(_01725_),
    .Y(_01731_)
  );
  AOI21X1 _08180_ (
    .A(_01720_),
    .B(_01731_),
    .C(_01717_),
    .Y(_01732_)
  );
  OAI21X1 _08181_ (
    .A(_01719_),
    .B(_01730_),
    .C(_01718_),
    .Y(_01733_)
  );
  XNOR2X1 _08182_ (
    .A(_01720_),
    .B(_01730_),
    .Y(_01734_)
  );
  XNOR2X1 _08183_ (
    .A(_01720_),
    .B(_01731_),
    .Y(_01735_)
  );
  XNOR2X1 _08184_ (
    .A(_01726_),
    .B(_01729_),
    .Y(_01736_)
  );
  NOR2X1 _08185_ (
    .A(_01714_),
    .B(_01736_),
    .Y(_01737_)
  );
  OR2X1 _08186_ (
    .A(_01714_),
    .B(_01736_),
    .Y(_01738_)
  );
  AOI21X1 _08187_ (
    .A(_01734_),
    .B(_01738_),
    .C(_01733_),
    .Y(_01739_)
  );
  OAI21X1 _08188_ (
    .A(_01735_),
    .B(_01737_),
    .C(_01732_),
    .Y(_01740_)
  );
  NOR2X1 _08189_ (
    .A(_01714_),
    .B(_01739_),
    .Y(_01741_)
  );
  XNOR2X1 _08190_ (
    .A(_01714_),
    .B(_01740_),
    .Y(_01742_)
  );
  NAND2X1 _08191_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01711_),
    .Y(_01743_)
  );
  NAND2X1 _08192_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01701_),
    .Y(_01744_)
  );
  AOI21X1 _08193_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_0_ ),
    .C(_01659_),
    .Y(_01745_)
  );
  OAI21X1 _08194_ (
    .A(_01413_),
    .B(_01704_),
    .C(_01745_),
    .Y(_01746_)
  );
  AOI22X1 _08195_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_9_ ),
    .C(_01453_),
    .D(_01700_),
    .Y(_01747_)
  );
  NAND3X1 _08196_ (
    .A(_01743_),
    .B(_01744_),
    .C(_01747_),
    .Y(_01748_)
  );
  OAI21X1 _08197_ (
    .A(_01746_),
    .B(_01748_),
    .C(_01424_),
    .Y(_01749_)
  );
  AOI22X1 _08198_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01742_),
    .C(_01749_),
    .D(_01542_),
    .Y(_01750_)
  );
  INVX1 _08199_ (
    .A(_01750_),
    .Y(_01751_)
  );
  OAI21X1 _08200_ (
    .A(_01708_),
    .B(_01710_),
    .C(_01751_),
    .Y(execution_unit_0.alu_0.alu_out_9_ )
  );
  NOR2X1 _08201_ (
    .A(_01678_),
    .B(_01704_),
    .Y(_01752_)
  );
  NOR2X1 _08202_ (
    .A(_01703_),
    .B(_01752_),
    .Y(_01753_)
  );
  OAI21X1 _08203_ (
    .A(_01681_),
    .B(_01705_),
    .C(_01753_),
    .Y(_01754_)
  );
  NAND2X1 _08204_ (
    .A(_01438_),
    .B(_01722_),
    .Y(_01755_)
  );
  NAND2X1 _08205_ (
    .A(_01438_),
    .B(_01724_),
    .Y(_01756_)
  );
  AOI22X1 _08206_ (
    .A(_01438_),
    .B(_01724_),
    .C(_01755_),
    .D(_01723_),
    .Y(_01757_)
  );
  NAND2X1 _08207_ (
    .A(_01754_),
    .B(_01757_),
    .Y(_01758_)
  );
  XNOR2X1 _08208_ (
    .A(_01754_),
    .B(_01757_),
    .Y(_01759_)
  );
  INVX1 _08209_ (
    .A(_01759_),
    .Y(dbg_0.UNUSED_eu_mab_10_ )
  );
  NAND2X1 _08210_ (
    .A(_01709_),
    .B(_01759_),
    .Y(_01760_)
  );
  OR2X1 _08211_ (
    .A(_01709_),
    .B(_01759_),
    .Y(_01761_)
  );
  NAND2X1 _08212_ (
    .A(_01760_),
    .B(_01761_),
    .Y(_01762_)
  );
  AOI21X1 _08213_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_1_ ),
    .C(_01659_),
    .Y(_01763_)
  );
  AOI22X1 _08214_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_10_ ),
    .C(_01453_),
    .D(_01722_),
    .Y(_01764_)
  );
  OAI21X1 _08215_ (
    .A(_01414_),
    .B(_01725_),
    .C(_01764_),
    .Y(_01765_)
  );
  OAI21X1 _08216_ (
    .A(_01413_),
    .B(_01728_),
    .C(_01763_),
    .Y(_01766_)
  );
  NOR2X1 _08217_ (
    .A(_01765_),
    .B(_01766_),
    .Y(_01767_)
  );
  AOI21X1 _08218_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01729_),
    .C(_01425_),
    .Y(_01768_)
  );
  NAND2X1 _08219_ (
    .A(_01767_),
    .B(_01768_),
    .Y(_01769_)
  );
  OAI21X1 _08220_ (
    .A(_01417_),
    .B(_01425_),
    .C(_01769_),
    .Y(_01770_)
  );
  AOI21X1 _08221_ (
    .A(_01736_),
    .B(_01741_),
    .C(_01417_),
    .Y(_01771_)
  );
  OAI21X1 _08222_ (
    .A(_01736_),
    .B(_01741_),
    .C(_01771_),
    .Y(_01772_)
  );
  AOI22X1 _08223_ (
    .A(_01425_),
    .B(_01762_),
    .C(_01770_),
    .D(_01772_),
    .Y(execution_unit_0.alu_0.alu_out_10_ )
  );
  OAI21X1 _08224_ (
    .A(_01439_),
    .B(_01725_),
    .C(_01758_),
    .Y(_01773_)
  );
  NOR2X1 _08225_ (
    .A(_01439_),
    .B(_01718_),
    .Y(_01774_)
  );
  AOI22X1 _08226_ (
    .A(execution_unit_0.alu_0.op_dst_11_ ),
    .B(_01673_),
    .C(_01716_),
    .D(_01438_),
    .Y(_01775_)
  );
  NOR2X1 _08227_ (
    .A(_01774_),
    .B(_01775_),
    .Y(_01776_)
  );
  XNOR2X1 _08228_ (
    .A(_01773_),
    .B(_01776_),
    .Y(_01777_)
  );
  INVX1 _08229_ (
    .A(_01777_),
    .Y(dbg_0.UNUSED_eu_mab_11_ )
  );
  NOR2X1 _08230_ (
    .A(_01761_),
    .B(_01777_),
    .Y(_01778_)
  );
  XNOR2X1 _08231_ (
    .A(_01761_),
    .B(_01777_),
    .Y(_01779_)
  );
  AOI21X1 _08232_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_2_ ),
    .C(_01659_),
    .Y(_01780_)
  );
  AOI22X1 _08233_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_11_ ),
    .C(_01453_),
    .D(_01716_),
    .Y(_01781_)
  );
  OAI21X1 _08234_ (
    .A(_01414_),
    .B(_01718_),
    .C(_01781_),
    .Y(_01782_)
  );
  OAI21X1 _08235_ (
    .A(_01413_),
    .B(_01719_),
    .C(_01780_),
    .Y(_01783_)
  );
  NOR2X1 _08236_ (
    .A(_01782_),
    .B(_01783_),
    .Y(_01784_)
  );
  AOI21X1 _08237_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01720_),
    .C(_01425_),
    .Y(_01785_)
  );
  NAND2X1 _08238_ (
    .A(_01784_),
    .B(_01785_),
    .Y(_01786_)
  );
  OAI21X1 _08239_ (
    .A(_01732_),
    .B(_01737_),
    .C(_01735_),
    .Y(_01787_)
  );
  AOI21X1 _08240_ (
    .A(_01734_),
    .B(_01738_),
    .C(_01417_),
    .Y(_01788_)
  );
  AOI22X1 _08241_ (
    .A(_01542_),
    .B(_01786_),
    .C(_01787_),
    .D(_01788_),
    .Y(_01789_)
  );
  AOI21X1 _08242_ (
    .A(_01425_),
    .B(_01779_),
    .C(_01789_),
    .Y(execution_unit_0.alu_0.alu_out_11_ )
  );
  AOI21X1 _08243_ (
    .A(_01756_),
    .B(_01758_),
    .C(_01775_),
    .Y(_01790_)
  );
  OR2X1 _08244_ (
    .A(_01774_),
    .B(_01790_),
    .Y(_01791_)
  );
  OAI21X1 _08245_ (
    .A(execution_unit_0.alu_0.alu_shift_11_ ),
    .B(_01426_),
    .C(_01673_),
    .Y(_01792_)
  );
  AOI21X1 _08246_ (
    .A(execution_unit_0.alu_0.alu_shift_11_ ),
    .B(_01426_),
    .C(_01792_),
    .Y(_01793_)
  );
  AND2X1 _08247_ (
    .A(execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01793_),
    .Y(_01794_)
  );
  NAND2X1 _08248_ (
    .A(execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01793_),
    .Y(_01795_)
  );
  AOI22X1 _08249_ (
    .A(execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01673_),
    .C(_01793_),
    .D(_01438_),
    .Y(_01796_)
  );
  AOI21X1 _08250_ (
    .A(_01438_),
    .B(_01794_),
    .C(_01796_),
    .Y(_01797_)
  );
  XOR2X1 _08251_ (
    .A(_01791_),
    .B(_01797_),
    .Y(dbg_0.UNUSED_eu_mab_12_ )
  );
  AND2X1 _08252_ (
    .A(_01778_),
    .B(dbg_0.UNUSED_eu_mab_12_ ),
    .Y(_01798_)
  );
  OAI21X1 _08253_ (
    .A(_01778_),
    .B(dbg_0.UNUSED_eu_mab_12_ ),
    .C(_01425_),
    .Y(_01799_)
  );
  OR2X1 _08254_ (
    .A(_01798_),
    .B(_01799_),
    .Y(_01800_)
  );
  AOI21X1 _08255_ (
    .A(execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01673_),
    .C(_01793_),
    .Y(_01801_)
  );
  NOR2X1 _08256_ (
    .A(_01794_),
    .B(_01801_),
    .Y(_01802_)
  );
  INVX1 _08257_ (
    .A(_01802_),
    .Y(_01803_)
  );
  NOR3X1 _08258_ (
    .A(_01732_),
    .B(_01735_),
    .C(_01737_),
    .Y(_01804_)
  );
  NAND3X1 _08259_ (
    .A(_01733_),
    .B(_01734_),
    .C(_01738_),
    .Y(_01805_)
  );
  NOR3X1 _08260_ (
    .A(_01739_),
    .B(_01803_),
    .C(_01804_),
    .Y(_01806_)
  );
  NAND3X1 _08261_ (
    .A(_01740_),
    .B(_01802_),
    .C(_01805_),
    .Y(_01807_)
  );
  OAI21X1 _08262_ (
    .A(_01739_),
    .B(_01804_),
    .C(_01803_),
    .Y(_01808_)
  );
  AND2X1 _08263_ (
    .A(_01807_),
    .B(_01808_),
    .Y(_01809_)
  );
  NAND2X1 _08264_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01802_),
    .Y(_01810_)
  );
  NAND2X1 _08265_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01794_),
    .Y(_01811_)
  );
  AOI21X1 _08266_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_3_ ),
    .C(_01659_),
    .Y(_01812_)
  );
  OAI21X1 _08267_ (
    .A(_01413_),
    .B(_01801_),
    .C(_01812_),
    .Y(_01813_)
  );
  AOI22X1 _08268_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_12_ ),
    .C(_01453_),
    .D(_01793_),
    .Y(_01814_)
  );
  NAND3X1 _08269_ (
    .A(_01810_),
    .B(_01811_),
    .C(_01814_),
    .Y(_01815_)
  );
  OAI21X1 _08270_ (
    .A(_01813_),
    .B(_01815_),
    .C(_01424_),
    .Y(_01816_)
  );
  OAI21X1 _08271_ (
    .A(_01417_),
    .B(_01425_),
    .C(_01816_),
    .Y(_01817_)
  );
  OAI21X1 _08272_ (
    .A(_01417_),
    .B(_01809_),
    .C(_01817_),
    .Y(_01818_)
  );
  OAI21X1 _08273_ (
    .A(_01798_),
    .B(_01799_),
    .C(_01818_),
    .Y(execution_unit_0.alu_0.alu_out_12_ )
  );
  XNOR2X1 _08274_ (
    .A(execution_unit_0.alu_0.alu_shift_12_ ),
    .B(_01426_),
    .Y(_01819_)
  );
  NOR2X1 _08275_ (
    .A(_01672_),
    .B(_01819_),
    .Y(_01820_)
  );
  AND2X1 _08276_ (
    .A(execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01820_),
    .Y(_01821_)
  );
  NAND2X1 _08277_ (
    .A(execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01820_),
    .Y(_01822_)
  );
  AOI21X1 _08278_ (
    .A(execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01673_),
    .C(_01820_),
    .Y(_01823_)
  );
  AOI22X1 _08279_ (
    .A(execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01673_),
    .C(_01820_),
    .D(_01438_),
    .Y(_01824_)
  );
  AOI21X1 _08280_ (
    .A(_01438_),
    .B(_01821_),
    .C(_01824_),
    .Y(_01825_)
  );
  AOI22X1 _08281_ (
    .A(_01438_),
    .B(_01794_),
    .C(_01797_),
    .D(_01791_),
    .Y(_01826_)
  );
  XNOR2X1 _08282_ (
    .A(_01825_),
    .B(_01826_),
    .Y(dbg_0.UNUSED_eu_mab_13_ )
  );
  NOR2X1 _08283_ (
    .A(_01798_),
    .B(dbg_0.UNUSED_eu_mab_13_ ),
    .Y(_01827_)
  );
  NAND2X1 _08284_ (
    .A(_01798_),
    .B(dbg_0.UNUSED_eu_mab_13_ ),
    .Y(_01828_)
  );
  OAI21X1 _08285_ (
    .A(execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01423_),
    .C(_01828_),
    .Y(_01829_)
  );
  NOR2X1 _08286_ (
    .A(_01827_),
    .B(_01829_),
    .Y(_01830_)
  );
  NOR2X1 _08287_ (
    .A(_01821_),
    .B(_01823_),
    .Y(_01831_)
  );
  INVX1 _08288_ (
    .A(_01831_),
    .Y(_01832_)
  );
  NAND2X1 _08289_ (
    .A(_01795_),
    .B(_01807_),
    .Y(_01833_)
  );
  AOI21X1 _08290_ (
    .A(_01795_),
    .B(_01807_),
    .C(_01832_),
    .Y(_01834_)
  );
  OAI21X1 _08291_ (
    .A(_01794_),
    .B(_01806_),
    .C(_01831_),
    .Y(_01835_)
  );
  XNOR2X1 _08292_ (
    .A(_01832_),
    .B(_01833_),
    .Y(_01836_)
  );
  XNOR2X1 _08293_ (
    .A(_01831_),
    .B(_01833_),
    .Y(_01837_)
  );
  XNOR2X1 _08294_ (
    .A(execution_unit_0.alu_0.alu_shift_14_ ),
    .B(_01426_),
    .Y(_01838_)
  );
  NOR2X1 _08295_ (
    .A(_01672_),
    .B(_01838_),
    .Y(_01839_)
  );
  INVX1 _08296_ (
    .A(_01839_),
    .Y(_01840_)
  );
  NOR2X1 _08297_ (
    .A(_01422_),
    .B(_01840_),
    .Y(_01841_)
  );
  NAND2X1 _08298_ (
    .A(execution_unit_0.alu_0.op_dst_15_ ),
    .B(_01839_),
    .Y(_01842_)
  );
  OAI21X1 _08299_ (
    .A(_01422_),
    .B(_01672_),
    .C(_01840_),
    .Y(_01843_)
  );
  XNOR2X1 _08300_ (
    .A(execution_unit_0.alu_0.alu_shift_13_ ),
    .B(_01426_),
    .Y(_01844_)
  );
  NOR2X1 _08301_ (
    .A(_01672_),
    .B(_01844_),
    .Y(_01845_)
  );
  OAI21X1 _08302_ (
    .A(_01957_),
    .B(_01421_),
    .C(execution_unit_0.alu_0.op_dst_14_ ),
    .Y(_01846_)
  );
  NOR2X1 _08303_ (
    .A(_01844_),
    .B(_01846_),
    .Y(_01847_)
  );
  NAND2X1 _08304_ (
    .A(execution_unit_0.alu_0.op_dst_14_ ),
    .B(_01845_),
    .Y(_01848_)
  );
  OAI21X1 _08305_ (
    .A(_01672_),
    .B(_01844_),
    .C(_01846_),
    .Y(_01849_)
  );
  AND2X1 _08306_ (
    .A(_01848_),
    .B(_01849_),
    .Y(_01850_)
  );
  OAI21X1 _08307_ (
    .A(_01844_),
    .B(_01846_),
    .C(_01849_),
    .Y(_01851_)
  );
  AOI21X1 _08308_ (
    .A(_01822_),
    .B(_01835_),
    .C(_01851_),
    .Y(_01852_)
  );
  OAI21X1 _08309_ (
    .A(_01821_),
    .B(_01834_),
    .C(_01850_),
    .Y(_01853_)
  );
  OAI21X1 _08310_ (
    .A(_01847_),
    .B(_01852_),
    .C(_01843_),
    .Y(_01854_)
  );
  AND2X1 _08311_ (
    .A(_01842_),
    .B(_01854_),
    .Y(_01855_)
  );
  OAI21X1 _08312_ (
    .A(_01422_),
    .B(_01840_),
    .C(_01854_),
    .Y(_01856_)
  );
  NOR3X1 _08313_ (
    .A(_01821_),
    .B(_01834_),
    .C(_01850_),
    .Y(_01857_)
  );
  NAND3X1 _08314_ (
    .A(_01822_),
    .B(_01835_),
    .C(_01851_),
    .Y(_01858_)
  );
  NAND2X1 _08315_ (
    .A(_01853_),
    .B(_01858_),
    .Y(_01859_)
  );
  AOI21X1 _08316_ (
    .A(_01853_),
    .B(_01858_),
    .C(_01836_),
    .Y(_01860_)
  );
  OAI21X1 _08317_ (
    .A(_01852_),
    .B(_01857_),
    .C(_01837_),
    .Y(_01861_)
  );
  AND2X1 _08318_ (
    .A(_01842_),
    .B(_01843_),
    .Y(_01862_)
  );
  OAI21X1 _08319_ (
    .A(_01422_),
    .B(_01840_),
    .C(_01843_),
    .Y(_01863_)
  );
  OAI21X1 _08320_ (
    .A(_01847_),
    .B(_01852_),
    .C(_01863_),
    .Y(_01864_)
  );
  NAND3X1 _08321_ (
    .A(_01848_),
    .B(_01853_),
    .C(_01862_),
    .Y(_01865_)
  );
  NAND3X1 _08322_ (
    .A(_01848_),
    .B(_01853_),
    .C(_01863_),
    .Y(_01866_)
  );
  OAI21X1 _08323_ (
    .A(_01847_),
    .B(_01852_),
    .C(_01862_),
    .Y(_01867_)
  );
  NAND2X1 _08324_ (
    .A(_01866_),
    .B(_01867_),
    .Y(_01868_)
  );
  AOI21X1 _08325_ (
    .A(_01864_),
    .B(_01865_),
    .C(_01860_),
    .Y(_01869_)
  );
  NAND3X1 _08326_ (
    .A(_01861_),
    .B(_01866_),
    .C(_01867_),
    .Y(_01870_)
  );
  AOI21X1 _08327_ (
    .A(_01855_),
    .B(_01870_),
    .C(_01836_),
    .Y(_01871_)
  );
  OAI21X1 _08328_ (
    .A(_01856_),
    .B(_01869_),
    .C(_01837_),
    .Y(_01872_)
  );
  NAND3X1 _08329_ (
    .A(_01836_),
    .B(_01855_),
    .C(_01868_),
    .Y(_01873_)
  );
  NAND3X1 _08330_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01872_),
    .C(_01873_),
    .Y(_01874_)
  );
  NAND2X1 _08331_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01831_),
    .Y(_01875_)
  );
  NAND2X1 _08332_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01821_),
    .Y(_01876_)
  );
  AOI21X1 _08333_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_4_ ),
    .C(_01659_),
    .Y(_01877_)
  );
  OAI21X1 _08334_ (
    .A(_01413_),
    .B(_01823_),
    .C(_01877_),
    .Y(_01878_)
  );
  AOI22X1 _08335_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_13_ ),
    .C(_01453_),
    .D(_01820_),
    .Y(_01879_)
  );
  NAND3X1 _08336_ (
    .A(_01875_),
    .B(_01876_),
    .C(_01879_),
    .Y(_01880_)
  );
  OAI21X1 _08337_ (
    .A(_01878_),
    .B(_01880_),
    .C(_01424_),
    .Y(_01881_)
  );
  OAI21X1 _08338_ (
    .A(_01417_),
    .B(_01425_),
    .C(_01881_),
    .Y(_01882_)
  );
  AOI21X1 _08339_ (
    .A(_01874_),
    .B(_01882_),
    .C(_01830_),
    .Y(_01883_)
  );
  INVX1 _08340_ (
    .A(_01883_),
    .Y(execution_unit_0.alu_0.alu_out_13_ )
  );
  NAND2X1 _08341_ (
    .A(_01438_),
    .B(_01845_),
    .Y(_01884_)
  );
  AOI22X1 _08342_ (
    .A(_01438_),
    .B(_01847_),
    .C(_01884_),
    .D(_01846_),
    .Y(_01885_)
  );
  OAI22X1 _08343_ (
    .A(_01439_),
    .B(_01822_),
    .C(_01824_),
    .D(_01826_),
    .Y(_01886_)
  );
  NAND2X1 _08344_ (
    .A(_01885_),
    .B(_01886_),
    .Y(_01887_)
  );
  XNOR2X1 _08345_ (
    .A(_01885_),
    .B(_01886_),
    .Y(_01888_)
  );
  INVX1 _08346_ (
    .A(_01888_),
    .Y(dbg_0.UNUSED_eu_mab_14_ )
  );
  AOI21X1 _08347_ (
    .A(_01856_),
    .B(_01860_),
    .C(_01417_),
    .Y(_01889_)
  );
  OAI21X1 _08348_ (
    .A(_01859_),
    .B(_01871_),
    .C(_01889_),
    .Y(_01890_)
  );
  NAND2X1 _08349_ (
    .A(execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_01849_),
    .Y(_01891_)
  );
  AOI21X1 _08350_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_5_ ),
    .C(_01659_),
    .Y(_01892_)
  );
  AOI22X1 _08351_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_14_ ),
    .C(_01453_),
    .D(_01845_),
    .Y(_01893_)
  );
  OAI21X1 _08352_ (
    .A(_01414_),
    .B(_01848_),
    .C(_01893_),
    .Y(_01894_)
  );
  AOI21X1 _08353_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01850_),
    .C(_01894_),
    .Y(_01895_)
  );
  NAND3X1 _08354_ (
    .A(_01891_),
    .B(_01892_),
    .C(_01895_),
    .Y(_01896_)
  );
  OAI21X1 _08355_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01896_),
    .C(_01424_),
    .Y(_01897_)
  );
  INVX1 _08356_ (
    .A(_01897_),
    .Y(_01898_)
  );
  OR2X1 _08357_ (
    .A(_01828_),
    .B(_01888_),
    .Y(_01899_)
  );
  AOI21X1 _08358_ (
    .A(_01828_),
    .B(_01888_),
    .C(_01424_),
    .Y(_01900_)
  );
  AND2X1 _08359_ (
    .A(_01899_),
    .B(_01900_),
    .Y(_01901_)
  );
  AOI21X1 _08360_ (
    .A(_01890_),
    .B(_01898_),
    .C(_01901_),
    .Y(_01902_)
  );
  INVX1 _08361_ (
    .A(_01902_),
    .Y(execution_unit_0.alu_0.alu_out_14_ )
  );
  OAI21X1 _08362_ (
    .A(_01439_),
    .B(_01848_),
    .C(_01887_),
    .Y(_01903_)
  );
  AOI22X1 _08363_ (
    .A(execution_unit_0.alu_0.op_dst_15_ ),
    .B(_01673_),
    .C(_01839_),
    .D(_01438_),
    .Y(_01904_)
  );
  AOI21X1 _08364_ (
    .A(_01438_),
    .B(_01841_),
    .C(_01904_),
    .Y(_01905_)
  );
  NAND2X1 _08365_ (
    .A(_01903_),
    .B(_01905_),
    .Y(_01906_)
  );
  XNOR2X1 _08366_ (
    .A(_01903_),
    .B(_01905_),
    .Y(_01907_)
  );
  INVX1 _08367_ (
    .A(_01907_),
    .Y(dbg_0.UNUSED_eu_mab_15_ )
  );
  NOR2X1 _08368_ (
    .A(_01899_),
    .B(_01907_),
    .Y(_01908_)
  );
  AND2X1 _08369_ (
    .A(_01899_),
    .B(_01907_),
    .Y(_01909_)
  );
  OAI21X1 _08370_ (
    .A(_01908_),
    .B(_01909_),
    .C(_01425_),
    .Y(_01910_)
  );
  NAND2X1 _08371_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_6_ ),
    .Y(_01911_)
  );
  AOI22X1 _08372_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(_01655_),
    .C(_01839_),
    .D(_01453_),
    .Y(_01912_)
  );
  AOI21X1 _08373_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01841_),
    .C(_01659_),
    .Y(_01913_)
  );
  NAND2X1 _08374_ (
    .A(_01911_),
    .B(_01912_),
    .Y(_01914_)
  );
  AOI21X1 _08375_ (
    .A(execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_01843_),
    .C(_01914_),
    .Y(_01915_)
  );
  NAND2X1 _08376_ (
    .A(_01913_),
    .B(_01915_),
    .Y(_01916_)
  );
  OAI21X1 _08377_ (
    .A(_01412_),
    .B(_01863_),
    .C(_01424_),
    .Y(_01917_)
  );
  OAI21X1 _08378_ (
    .A(_01916_),
    .B(_01917_),
    .C(_01542_),
    .Y(_01918_)
  );
  AOI22X1 _08379_ (
    .A(_01856_),
    .B(_01861_),
    .C(_01866_),
    .D(_01867_),
    .Y(_01919_)
  );
  OAI21X1 _08380_ (
    .A(_01860_),
    .B(_01868_),
    .C(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01920_)
  );
  OAI21X1 _08381_ (
    .A(_01919_),
    .B(_01920_),
    .C(_01918_),
    .Y(_01921_)
  );
  NAND2X1 _08382_ (
    .A(_01910_),
    .B(_01921_),
    .Y(_01922_)
  );
  INVX1 _08383_ (
    .A(_01922_),
    .Y(execution_unit_0.alu_0.alu_out_15_ )
  );
  NAND2X1 _08384_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(execution_unit_0.alu_0.alu_out_7_ ),
    .Y(_01923_)
  );
  OAI21X1 _08385_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(_01922_),
    .C(_01923_),
    .Y(execution_unit_0.alu_0.N )
  );
  OR2X1 _08386_ (
    .A(execution_unit_0.alu_0.alu_out_8_ ),
    .B(execution_unit_0.alu_0.alu_out_11_ ),
    .Y(_01924_)
  );
  NOR3X1 _08387_ (
    .A(execution_unit_0.alu_0.alu_out_9_ ),
    .B(execution_unit_0.alu_0.alu_out_10_ ),
    .C(_01924_),
    .Y(_01925_)
  );
  NAND3X1 _08388_ (
    .A(_01800_),
    .B(_01818_),
    .C(_01925_),
    .Y(_01926_)
  );
  AOI21X1 _08389_ (
    .A(_01910_),
    .B(_01921_),
    .C(_01926_),
    .Y(_01927_)
  );
  NAND3X1 _08390_ (
    .A(_01883_),
    .B(_01902_),
    .C(_01927_),
    .Y(_01928_)
  );
  NOR2X1 _08391_ (
    .A(execution_unit_0.alu_0.alu_out_0_ ),
    .B(execution_unit_0.alu_0.alu_out_3_ ),
    .Y(_01929_)
  );
  NAND2X1 _08392_ (
    .A(_01516_),
    .B(_01929_),
    .Y(_01930_)
  );
  NOR2X1 _08393_ (
    .A(execution_unit_0.alu_0.alu_out_2_ ),
    .B(execution_unit_0.alu_0.alu_out_7_ ),
    .Y(_01931_)
  );
  NOR2X1 _08394_ (
    .A(execution_unit_0.alu_0.alu_out_4_ ),
    .B(_01930_),
    .Y(_01932_)
  );
  NAND2X1 _08395_ (
    .A(_01931_),
    .B(_01932_),
    .Y(_01933_)
  );
  OR2X1 _08396_ (
    .A(execution_unit_0.alu_0.alu_out_5_ ),
    .B(_01933_),
    .Y(_01934_)
  );
  OR2X1 _08397_ (
    .A(execution_unit_0.alu_0.alu_out_6_ ),
    .B(_01934_),
    .Y(_01935_)
  );
  AOI21X1 _08398_ (
    .A(_01421_),
    .B(_01928_),
    .C(_01935_),
    .Y(execution_unit_0.alu_0.Z )
  );
  NAND2X1 _08399_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(_01428_),
    .Y(_01936_)
  );
  OR2X1 _08400_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(execution_unit_0.alu_0.inst_alu_8_ ),
    .Y(_01937_)
  );
  AND2X1 _08401_ (
    .A(execution_unit_0.alu_0.Z ),
    .B(_01937_),
    .Y(_01938_)
  );
  OAI21X1 _08402_ (
    .A(_01439_),
    .B(_01842_),
    .C(_01906_),
    .Y(_01939_)
  );
  OAI21X1 _08403_ (
    .A(_01908_),
    .B(_01939_),
    .C(_01425_),
    .Y(_01940_)
  );
  AOI21X1 _08404_ (
    .A(_01855_),
    .B(_01870_),
    .C(_01542_),
    .Y(_01941_)
  );
  OAI21X1 _08405_ (
    .A(_01855_),
    .B(_01870_),
    .C(_01941_),
    .Y(_01942_)
  );
  AOI21X1 _08406_ (
    .A(_01940_),
    .B(_01942_),
    .C(execution_unit_0.alu_0.inst_bw ),
    .Y(_01943_)
  );
  AND2X1 _08407_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(execution_unit_0.alu_0.alu_out_8_ ),
    .Y(_01944_)
  );
  OR2X1 _08408_ (
    .A(_01943_),
    .B(_01944_),
    .Y(_01945_)
  );
  OAI21X1 _08409_ (
    .A(_01937_),
    .B(_01945_),
    .C(_01415_),
    .Y(_01946_)
  );
  OAI21X1 _08410_ (
    .A(_01938_),
    .B(_01946_),
    .C(_01936_),
    .Y(execution_unit_0.alu_0.alu_stat_0_ )
  );
  OAI21X1 _08411_ (
    .A(execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01604_),
    .C(execution_unit_0.alu_0.alu_out_7_ ),
    .Y(_01947_)
  );
  OAI21X1 _08412_ (
    .A(_01605_),
    .B(execution_unit_0.alu_0.alu_out_7_ ),
    .C(_01947_),
    .Y(_01948_)
  );
  NAND2X1 _08413_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(_01948_),
    .Y(_01949_)
  );
  NAND2X1 _08414_ (
    .A(_01841_),
    .B(_01922_),
    .Y(_01950_)
  );
  OAI21X1 _08415_ (
    .A(_01843_),
    .B(_01922_),
    .C(_01950_),
    .Y(_01951_)
  );
  OAI21X1 _08416_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(_01951_),
    .C(_01949_),
    .Y(_01952_)
  );
  AOI21X1 _08417_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(_01605_),
    .C(_01412_),
    .Y(_01953_)
  );
  OAI21X1 _08418_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(_01842_),
    .C(_01953_),
    .Y(_01954_)
  );
  NOR2X1 _08419_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.inst_alu_8_ ),
    .Y(_01955_)
  );
  NAND2X1 _08420_ (
    .A(_01954_),
    .B(_01955_),
    .Y(_01956_)
  );
  AOI21X1 _08421_ (
    .A(_01412_),
    .B(_01952_),
    .C(_01956_),
    .Y(execution_unit_0.alu_0.alu_stat_3_ )
  );
  AND2X1 _08422_ (
    .A(execution_unit_0.alu_0.exec_cycle ),
    .B(execution_unit_0.alu_0.inst_alu_9_ ),
    .Y(execution_unit_0.alu_0.alu_stat_wr_0_ )
  );
  INVX1 _08423_ (
    .A(execution_unit_0.reg_sr_clr ),
    .Y(_02980_)
  );
  INVX1 _08424_ (
    .A(execution_unit_0.inst_src_1_ ),
    .Y(_02981_)
  );
  INVX1 _08425_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .Y(_02982_)
  );
  INVX1 _08426_ (
    .A(execution_unit_0.register_file_0.r7_0_ ),
    .Y(_02983_)
  );
  INVX1 _08427_ (
    .A(execution_unit_0.alu_0.alu_out_0_ ),
    .Y(_02984_)
  );
  INVX1 _08428_ (
    .A(execution_unit_0.register_file_0.r1_1_ ),
    .Y(_02985_)
  );
  INVX1 _08429_ (
    .A(execution_unit_0.register_file_0.r4_1_ ),
    .Y(_02986_)
  );
  INVX1 _08430_ (
    .A(execution_unit_0.register_file_0.r7_1_ ),
    .Y(_02987_)
  );
  INVX1 _08431_ (
    .A(execution_unit_0.register_file_0.r10_1_ ),
    .Y(_02988_)
  );
  INVX1 _08432_ (
    .A(execution_unit_0.alu_0.alu_out_1_ ),
    .Y(_02989_)
  );
  INVX1 _08433_ (
    .A(execution_unit_0.register_file_0.r10_2_ ),
    .Y(_02990_)
  );
  INVX1 _08434_ (
    .A(execution_unit_0.alu_0.alu_out_2_ ),
    .Y(_02991_)
  );
  INVX1 _08435_ (
    .A(execution_unit_0.register_file_0.r1_3_ ),
    .Y(_02992_)
  );
  INVX1 _08436_ (
    .A(execution_unit_0.register_file_0.r7_3_ ),
    .Y(_02993_)
  );
  INVX1 _08437_ (
    .A(execution_unit_0.register_file_0.r13_3_ ),
    .Y(_02994_)
  );
  INVX1 _08438_ (
    .A(execution_unit_0.alu_0.alu_out_3_ ),
    .Y(_02995_)
  );
  INVX1 _08439_ (
    .A(execution_unit_0.register_file_0.r2_4_ ),
    .Y(_02996_)
  );
  INVX1 _08440_ (
    .A(execution_unit_0.register_file_0.r1_4_ ),
    .Y(_02997_)
  );
  INVX1 _08441_ (
    .A(execution_unit_0.alu_0.alu_out_4_ ),
    .Y(_02998_)
  );
  INVX1 _08442_ (
    .A(execution_unit_0.register_file_0.r1_5_ ),
    .Y(_02999_)
  );
  INVX1 _08443_ (
    .A(execution_unit_0.alu_0.alu_out_5_ ),
    .Y(_03000_)
  );
  INVX1 _08444_ (
    .A(execution_unit_0.register_file_0.r1_6_ ),
    .Y(_03001_)
  );
  INVX1 _08445_ (
    .A(execution_unit_0.alu_0.alu_out_6_ ),
    .Y(_03002_)
  );
  INVX1 _08446_ (
    .A(execution_unit_0.register_file_0.r1_7_ ),
    .Y(_03003_)
  );
  INVX1 _08447_ (
    .A(execution_unit_0.alu_0.alu_out_7_ ),
    .Y(_03004_)
  );
  INVX1 _08448_ (
    .A(execution_unit_0.register_file_0.r1_8_ ),
    .Y(_03005_)
  );
  INVX1 _08449_ (
    .A(execution_unit_0.register_file_0.r1_9_ ),
    .Y(_03006_)
  );
  INVX1 _08450_ (
    .A(execution_unit_0.register_file_0.r13_9_ ),
    .Y(_03007_)
  );
  INVX1 _08451_ (
    .A(execution_unit_0.register_file_0.r4_10_ ),
    .Y(_03008_)
  );
  INVX1 _08452_ (
    .A(execution_unit_0.register_file_0.r1_11_ ),
    .Y(_03009_)
  );
  INVX1 _08453_ (
    .A(execution_unit_0.register_file_0.r1_12_ ),
    .Y(_03010_)
  );
  INVX1 _08454_ (
    .A(execution_unit_0.register_file_0.r1_13_ ),
    .Y(_03011_)
  );
  INVX1 _08455_ (
    .A(execution_unit_0.register_file_0.r1_14_ ),
    .Y(_03012_)
  );
  INVX1 _08456_ (
    .A(execution_unit_0.register_file_0.r10_14_ ),
    .Y(_03013_)
  );
  INVX1 _08457_ (
    .A(execution_unit_0.register_file_0.r13_15_ ),
    .Y(_03014_)
  );
  INVX1 _08458_ (
    .A(execution_unit_0.register_file_0.r1_15_ ),
    .Y(_03015_)
  );
  INVX1 _08459_ (
    .A(execution_unit_0.reg_sp_wr ),
    .Y(_03016_)
  );
  INVX1 _08460_ (
    .A(execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .Y(_03017_)
  );
  INVX1 _08461_ (
    .A(execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .Y(_03018_)
  );
  INVX1 _08462_ (
    .A(execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .Y(_03019_)
  );
  INVX1 _08463_ (
    .A(execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .Y(_03020_)
  );
  INVX1 _08464_ (
    .A(_00162_),
    .Y(_02190_)
  );
  AND2X1 _08465_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_6_ ),
    .Y(_03021_)
  );
  NAND3X1 _08466_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_6_ ),
    .C(execution_unit_0.register_file_0.r6_0_ ),
    .Y(_03022_)
  );
  AND2X1 _08467_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_11_ ),
    .Y(_03023_)
  );
  NAND3X1 _08468_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_11_ ),
    .C(execution_unit_0.register_file_0.r11_0_ ),
    .Y(_03024_)
  );
  AND2X1 _08469_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_9_ ),
    .Y(_03025_)
  );
  NAND3X1 _08470_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_9_ ),
    .C(execution_unit_0.register_file_0.r9_0_ ),
    .Y(_03026_)
  );
  AND2X1 _08471_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_3_ ),
    .Y(_03027_)
  );
  AND2X1 _08472_ (
    .A(execution_unit_0.register_file_0.r3_0_ ),
    .B(_03027_),
    .Y(_03028_)
  );
  AND2X1 _08473_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_12_ ),
    .Y(_03029_)
  );
  NAND3X1 _08474_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_12_ ),
    .C(execution_unit_0.register_file_0.r12_0_ ),
    .Y(_03030_)
  );
  NOR2X1 _08475_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(_02981_),
    .Y(_03031_)
  );
  NAND3X1 _08476_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_1_ ),
    .C(execution_unit_0.register_file_0.r1_0_ ),
    .Y(_03032_)
  );
  OR2X1 _08477_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(execution_unit_0.inst_src_2_ ),
    .Y(_03033_)
  );
  AND2X1 _08478_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_8_ ),
    .Y(_03034_)
  );
  NAND3X1 _08479_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_8_ ),
    .C(execution_unit_0.register_file_0.r8_0_ ),
    .Y(_03035_)
  );
  AND2X1 _08480_ (
    .A(execution_unit_0.inst_src_14_ ),
    .B(_02980_),
    .Y(_03036_)
  );
  NAND3X1 _08481_ (
    .A(execution_unit_0.inst_src_14_ ),
    .B(_02980_),
    .C(execution_unit_0.register_file_0.r14_0_ ),
    .Y(_03037_)
  );
  AND2X1 _08482_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_13_ ),
    .Y(_03038_)
  );
  NAND2X1 _08483_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_13_ ),
    .Y(_03039_)
  );
  NAND3X1 _08484_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_13_ ),
    .C(execution_unit_0.register_file_0.r13_0_ ),
    .Y(_03040_)
  );
  AND2X1 _08485_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_4_ ),
    .Y(_03041_)
  );
  NAND2X1 _08486_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_4_ ),
    .Y(_03042_)
  );
  NAND3X1 _08487_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_4_ ),
    .C(execution_unit_0.register_file_0.r4_0_ ),
    .Y(_03043_)
  );
  AND2X1 _08488_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_10_ ),
    .Y(_03044_)
  );
  NAND2X1 _08489_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_10_ ),
    .Y(_03045_)
  );
  NAND3X1 _08490_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_10_ ),
    .C(execution_unit_0.register_file_0.r10_0_ ),
    .Y(_03046_)
  );
  AND2X1 _08491_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_7_ ),
    .Y(_03047_)
  );
  NAND2X1 _08492_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_7_ ),
    .Y(_03048_)
  );
  AND2X1 _08493_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_0_ ),
    .Y(_03049_)
  );
  NAND3X1 _08494_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_0_ ),
    .C(dbg_0.UNUSED_pc_0_ ),
    .Y(_03050_)
  );
  OAI21X1 _08495_ (
    .A(_02983_),
    .B(_03048_),
    .C(_03050_),
    .Y(_03051_)
  );
  AND2X1 _08496_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_15_ ),
    .Y(_03052_)
  );
  NAND3X1 _08497_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_15_ ),
    .C(execution_unit_0.register_file_0.r15_0_ ),
    .Y(_03053_)
  );
  AND2X1 _08498_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_5_ ),
    .Y(_03054_)
  );
  NAND3X1 _08499_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_5_ ),
    .C(execution_unit_0.register_file_0.r5_0_ ),
    .Y(_03055_)
  );
  NAND3X1 _08500_ (
    .A(_03030_),
    .B(_03032_),
    .C(_03037_),
    .Y(_03056_)
  );
  NAND3X1 _08501_ (
    .A(_03022_),
    .B(_03024_),
    .C(_03040_),
    .Y(_03057_)
  );
  NOR2X1 _08502_ (
    .A(_03056_),
    .B(_03057_),
    .Y(_03058_)
  );
  NAND3X1 _08503_ (
    .A(_03026_),
    .B(_03053_),
    .C(_03055_),
    .Y(_03059_)
  );
  NOR3X1 _08504_ (
    .A(_03028_),
    .B(_03051_),
    .C(_03059_),
    .Y(_03060_)
  );
  NAND3X1 _08505_ (
    .A(_03035_),
    .B(_03043_),
    .C(_03046_),
    .Y(_03061_)
  );
  AOI21X1 _08506_ (
    .A(execution_unit_0.alu_0.status_0_ ),
    .B(_03033_),
    .C(_03061_),
    .Y(_03062_)
  );
  NAND3X1 _08507_ (
    .A(_03058_),
    .B(_03060_),
    .C(_03062_),
    .Y(execution_unit_0.reg_src_0_ )
  );
  AND2X1 _08508_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.reg_dest_wr ),
    .Y(_03063_)
  );
  NAND2X1 _08509_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.reg_dest_wr ),
    .Y(_03064_)
  );
  AND2X1 _08510_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03036_),
    .Y(_03065_)
  );
  NAND2X1 _08511_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03036_),
    .Y(_03066_)
  );
  OAI21X1 _08512_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(_02981_),
    .C(execution_unit_0.alu_0.inst_bw ),
    .Y(_03067_)
  );
  NOR2X1 _08513_ (
    .A(execution_unit_0.reg_src_0_ ),
    .B(_03067_),
    .Y(_03068_)
  );
  XOR2X1 _08514_ (
    .A(execution_unit_0.reg_src_0_ ),
    .B(_03067_),
    .Y(_03069_)
  );
  AOI21X1 _08515_ (
    .A(_03065_),
    .B(_03069_),
    .C(_03063_),
    .Y(_03070_)
  );
  OAI21X1 _08516_ (
    .A(execution_unit_0.register_file_0.r14_0_ ),
    .B(_03065_),
    .C(_03070_),
    .Y(_03071_)
  );
  OAI21X1 _08517_ (
    .A(_02984_),
    .B(_03064_),
    .C(_03071_),
    .Y(_02022_)
  );
  NAND3X1 _08518_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_0_ ),
    .C(dbg_0.UNUSED_pc_1_ ),
    .Y(_03072_)
  );
  NAND3X1 _08519_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_3_ ),
    .C(execution_unit_0.register_file_0.r3_1_ ),
    .Y(_03073_)
  );
  NAND3X1 _08520_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_1_ ),
    .C(execution_unit_0.register_file_0.r1_1_ ),
    .Y(_03074_)
  );
  NAND3X1 _08521_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_8_ ),
    .C(execution_unit_0.register_file_0.r8_1_ ),
    .Y(_03075_)
  );
  OAI21X1 _08522_ (
    .A(_02986_),
    .B(_03042_),
    .C(_03075_),
    .Y(_03076_)
  );
  AND2X1 _08523_ (
    .A(execution_unit_0.register_file_0.r14_1_ ),
    .B(_03036_),
    .Y(_03077_)
  );
  NAND2X1 _08524_ (
    .A(execution_unit_0.register_file_0.r12_1_ ),
    .B(_03029_),
    .Y(_03078_)
  );
  NAND3X1 _08525_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_13_ ),
    .C(execution_unit_0.register_file_0.r13_1_ ),
    .Y(_03079_)
  );
  NAND3X1 _08526_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_15_ ),
    .C(execution_unit_0.register_file_0.r15_1_ ),
    .Y(_03080_)
  );
  OAI21X1 _08527_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(execution_unit_0.inst_src_2_ ),
    .C(execution_unit_0.alu_0.status_1_ ),
    .Y(_03081_)
  );
  NAND3X1 _08528_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_11_ ),
    .C(execution_unit_0.register_file_0.r11_1_ ),
    .Y(_03082_)
  );
  NAND3X1 _08529_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_5_ ),
    .C(execution_unit_0.register_file_0.r5_1_ ),
    .Y(_03083_)
  );
  NAND3X1 _08530_ (
    .A(_03079_),
    .B(_03080_),
    .C(_03082_),
    .Y(_03084_)
  );
  NAND3X1 _08531_ (
    .A(_03073_),
    .B(_03081_),
    .C(_03083_),
    .Y(_03085_)
  );
  OAI21X1 _08532_ (
    .A(_02987_),
    .B(_03048_),
    .C(_03074_),
    .Y(_03086_)
  );
  NOR3X1 _08533_ (
    .A(_03084_),
    .B(_03085_),
    .C(_03086_),
    .Y(_03087_)
  );
  AOI22X1 _08534_ (
    .A(execution_unit_0.register_file_0.r6_1_ ),
    .B(_03021_),
    .C(_03025_),
    .D(execution_unit_0.register_file_0.r9_1_ ),
    .Y(_03088_)
  );
  AND2X1 _08535_ (
    .A(_03078_),
    .B(_03088_),
    .Y(_03089_)
  );
  OAI21X1 _08536_ (
    .A(_02988_),
    .B(_03045_),
    .C(_03072_),
    .Y(_03090_)
  );
  NOR3X1 _08537_ (
    .A(_03076_),
    .B(_03077_),
    .C(_03090_),
    .Y(_03091_)
  );
  NAND3X1 _08538_ (
    .A(_03087_),
    .B(_03089_),
    .C(_03091_),
    .Y(execution_unit_0.reg_src_1_ )
  );
  OAI21X1 _08539_ (
    .A(execution_unit_0.reg_src_0_ ),
    .B(_03067_),
    .C(execution_unit_0.reg_src_1_ ),
    .Y(_03092_)
  );
  XNOR2X1 _08540_ (
    .A(_03068_),
    .B(execution_unit_0.reg_src_1_ ),
    .Y(_03093_)
  );
  NOR2X1 _08541_ (
    .A(execution_unit_0.register_file_0.r14_1_ ),
    .B(_03065_),
    .Y(_03094_)
  );
  OAI21X1 _08542_ (
    .A(_03066_),
    .B(_03093_),
    .C(_03064_),
    .Y(_03095_)
  );
  OAI22X1 _08543_ (
    .A(_02989_),
    .B(_03064_),
    .C(_03094_),
    .D(_03095_),
    .Y(_02029_)
  );
  NAND2X1 _08544_ (
    .A(execution_unit_0.register_file_0.r9_2_ ),
    .B(_03025_),
    .Y(_03096_)
  );
  AOI22X1 _08545_ (
    .A(execution_unit_0.register_file_0.r13_2_ ),
    .B(_03038_),
    .C(_03047_),
    .D(execution_unit_0.register_file_0.r7_2_ ),
    .Y(_03097_)
  );
  AOI22X1 _08546_ (
    .A(execution_unit_0.register_file_0.r4_2_ ),
    .B(_03041_),
    .C(_03052_),
    .D(execution_unit_0.register_file_0.r15_2_ ),
    .Y(_03098_)
  );
  AOI22X1 _08547_ (
    .A(execution_unit_0.register_file_0.r11_2_ ),
    .B(_03023_),
    .C(_03034_),
    .D(execution_unit_0.register_file_0.r8_2_ ),
    .Y(_03099_)
  );
  AOI22X1 _08548_ (
    .A(execution_unit_0.register_file_0.r12_2_ ),
    .B(_03029_),
    .C(_03036_),
    .D(execution_unit_0.register_file_0.r14_2_ ),
    .Y(_03100_)
  );
  NAND2X1 _08549_ (
    .A(_03099_),
    .B(_03100_),
    .Y(_03101_)
  );
  NAND2X1 _08550_ (
    .A(_03096_),
    .B(_03097_),
    .Y(_03102_)
  );
  AOI22X1 _08551_ (
    .A(execution_unit_0.register_file_0.r3_2_ ),
    .B(_03027_),
    .C(_03049_),
    .D(dbg_0.UNUSED_pc_2_ ),
    .Y(_03103_)
  );
  OAI21X1 _08552_ (
    .A(_02990_),
    .B(_03045_),
    .C(_03103_),
    .Y(_03104_)
  );
  NOR2X1 _08553_ (
    .A(_03102_),
    .B(_03104_),
    .Y(_03105_)
  );
  AOI22X1 _08554_ (
    .A(execution_unit_0.alu_0.status_2_ ),
    .B(_03033_),
    .C(_03054_),
    .D(execution_unit_0.register_file_0.r5_2_ ),
    .Y(_03106_)
  );
  AOI22X1 _08555_ (
    .A(execution_unit_0.register_file_0.r6_2_ ),
    .B(_03021_),
    .C(_03031_),
    .D(execution_unit_0.register_file_0.r1_2_ ),
    .Y(_03107_)
  );
  NAND3X1 _08556_ (
    .A(_03098_),
    .B(_03106_),
    .C(_03107_),
    .Y(_03108_)
  );
  NOR2X1 _08557_ (
    .A(_03101_),
    .B(_03108_),
    .Y(_03109_)
  );
  AND2X1 _08558_ (
    .A(_03105_),
    .B(_03109_),
    .Y(_03110_)
  );
  INVX1 _08559_ (
    .A(_03110_),
    .Y(execution_unit_0.reg_src_2_ )
  );
  NOR2X1 _08560_ (
    .A(_03092_),
    .B(_03110_),
    .Y(_03111_)
  );
  XNOR2X1 _08561_ (
    .A(_03092_),
    .B(_03110_),
    .Y(_03112_)
  );
  AND2X1 _08562_ (
    .A(_03065_),
    .B(_03112_),
    .Y(_03113_)
  );
  OAI21X1 _08563_ (
    .A(execution_unit_0.register_file_0.r14_2_ ),
    .B(_03065_),
    .C(_03064_),
    .Y(_03114_)
  );
  OAI22X1 _08564_ (
    .A(_02991_),
    .B(_03064_),
    .C(_03113_),
    .D(_03114_),
    .Y(_02030_)
  );
  NAND2X1 _08565_ (
    .A(execution_unit_0.register_file_0.r5_3_ ),
    .B(_03054_),
    .Y(_03115_)
  );
  NAND3X1 _08566_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_9_ ),
    .C(execution_unit_0.register_file_0.r9_3_ ),
    .Y(_03116_)
  );
  NAND3X1 _08567_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_11_ ),
    .C(execution_unit_0.register_file_0.r11_3_ ),
    .Y(_03117_)
  );
  NAND2X1 _08568_ (
    .A(execution_unit_0.register_file_0.r6_3_ ),
    .B(_03021_),
    .Y(_03118_)
  );
  NAND3X1 _08569_ (
    .A(_02980_),
    .B(execution_unit_0.inst_src_12_ ),
    .C(execution_unit_0.register_file_0.r12_3_ ),
    .Y(_03119_)
  );
  NAND2X1 _08570_ (
    .A(execution_unit_0.register_file_0.r10_3_ ),
    .B(_03044_),
    .Y(_03120_)
  );
  AOI22X1 _08571_ (
    .A(execution_unit_0.register_file_0.r4_3_ ),
    .B(_03041_),
    .C(_03052_),
    .D(execution_unit_0.register_file_0.r15_3_ ),
    .Y(_03121_)
  );
  OAI22X1 _08572_ (
    .A(_02994_),
    .B(_03039_),
    .C(_03048_),
    .D(_02993_),
    .Y(_03122_)
  );
  NAND3X1 _08573_ (
    .A(_03116_),
    .B(_03117_),
    .C(_03119_),
    .Y(_03123_)
  );
  AOI21X1 _08574_ (
    .A(execution_unit_0.register_file_0.r8_3_ ),
    .B(_03034_),
    .C(_03123_),
    .Y(_03124_)
  );
  AOI21X1 _08575_ (
    .A(execution_unit_0.register_file_0.r14_3_ ),
    .B(_03036_),
    .C(_03122_),
    .Y(_03125_)
  );
  AOI22X1 _08576_ (
    .A(execution_unit_0.register_file_0.r3_3_ ),
    .B(_03027_),
    .C(_03049_),
    .D(dbg_0.UNUSED_pc_3_ ),
    .Y(_03126_)
  );
  AND2X1 _08577_ (
    .A(_03120_),
    .B(_03126_),
    .Y(_03127_)
  );
  NAND3X1 _08578_ (
    .A(_03124_),
    .B(_03125_),
    .C(_03127_),
    .Y(_03128_)
  );
  AOI22X1 _08579_ (
    .A(execution_unit_0.register_file_0.r1_3_ ),
    .B(_03031_),
    .C(_03033_),
    .D(execution_unit_0.gie ),
    .Y(_03129_)
  );
  AND2X1 _08580_ (
    .A(_03121_),
    .B(_03129_),
    .Y(_03130_)
  );
  NAND3X1 _08581_ (
    .A(_03115_),
    .B(_03118_),
    .C(_03130_),
    .Y(_03131_)
  );
  NOR2X1 _08582_ (
    .A(_03128_),
    .B(_03131_),
    .Y(_03132_)
  );
  INVX1 _08583_ (
    .A(_03132_),
    .Y(execution_unit_0.reg_src_3_ )
  );
  NOR3X1 _08584_ (
    .A(_03092_),
    .B(_03110_),
    .C(_03132_),
    .Y(_03133_)
  );
  NOR2X1 _08585_ (
    .A(_03111_),
    .B(execution_unit_0.reg_src_3_ ),
    .Y(_03134_)
  );
  NOR2X1 _08586_ (
    .A(_03133_),
    .B(_03134_),
    .Y(_03135_)
  );
  NOR2X1 _08587_ (
    .A(execution_unit_0.register_file_0.r14_3_ ),
    .B(_03065_),
    .Y(_03136_)
  );
  OAI21X1 _08588_ (
    .A(_03066_),
    .B(_03135_),
    .C(_03064_),
    .Y(_03137_)
  );
  OAI22X1 _08589_ (
    .A(_02995_),
    .B(_03064_),
    .C(_03136_),
    .D(_03137_),
    .Y(_02031_)
  );
  AOI22X1 _08590_ (
    .A(execution_unit_0.register_file_0.r4_4_ ),
    .B(_03041_),
    .C(_03049_),
    .D(dbg_0.UNUSED_pc_4_ ),
    .Y(_03138_)
  );
  AOI22X1 _08591_ (
    .A(execution_unit_0.register_file_0.r12_4_ ),
    .B(_03029_),
    .C(_03036_),
    .D(execution_unit_0.register_file_0.r14_4_ ),
    .Y(_03139_)
  );
  NAND2X1 _08592_ (
    .A(_03138_),
    .B(_03139_),
    .Y(_03140_)
  );
  AOI22X1 _08593_ (
    .A(execution_unit_0.register_file_0.r3_4_ ),
    .B(_03027_),
    .C(_03031_),
    .D(execution_unit_0.register_file_0.r1_4_ ),
    .Y(_03141_)
  );
  AOI22X1 _08594_ (
    .A(execution_unit_0.register_file_0.r9_4_ ),
    .B(_03025_),
    .C(_03054_),
    .D(execution_unit_0.register_file_0.r5_4_ ),
    .Y(_03142_)
  );
  NAND2X1 _08595_ (
    .A(_03141_),
    .B(_03142_),
    .Y(_03143_)
  );
  NOR2X1 _08596_ (
    .A(_03140_),
    .B(_03143_),
    .Y(_03144_)
  );
  AOI22X1 _08597_ (
    .A(execution_unit_0.register_file_0.r13_4_ ),
    .B(_03038_),
    .C(_03047_),
    .D(execution_unit_0.register_file_0.r7_4_ ),
    .Y(_03145_)
  );
  AOI22X1 _08598_ (
    .A(execution_unit_0.register_file_0.r6_4_ ),
    .B(_03021_),
    .C(_03034_),
    .D(execution_unit_0.register_file_0.r8_4_ ),
    .Y(_03146_)
  );
  NAND2X1 _08599_ (
    .A(_03145_),
    .B(_03146_),
    .Y(_03147_)
  );
  AOI22X1 _08600_ (
    .A(execution_unit_0.register_file_0.r2_4_ ),
    .B(_03033_),
    .C(_03052_),
    .D(execution_unit_0.register_file_0.r15_4_ ),
    .Y(_03148_)
  );
  AOI22X1 _08601_ (
    .A(execution_unit_0.register_file_0.r11_4_ ),
    .B(_03023_),
    .C(_03044_),
    .D(execution_unit_0.register_file_0.r10_4_ ),
    .Y(_03149_)
  );
  NAND2X1 _08602_ (
    .A(_03148_),
    .B(_03149_),
    .Y(_03150_)
  );
  NOR2X1 _08603_ (
    .A(_03147_),
    .B(_03150_),
    .Y(_03151_)
  );
  NAND2X1 _08604_ (
    .A(_03144_),
    .B(_03151_),
    .Y(execution_unit_0.reg_src_4_ )
  );
  NAND2X1 _08605_ (
    .A(_03133_),
    .B(execution_unit_0.reg_src_4_ ),
    .Y(_03152_)
  );
  XOR2X1 _08606_ (
    .A(_03133_),
    .B(execution_unit_0.reg_src_4_ ),
    .Y(_03153_)
  );
  NOR2X1 _08607_ (
    .A(execution_unit_0.register_file_0.r14_4_ ),
    .B(_03065_),
    .Y(_03154_)
  );
  OAI21X1 _08608_ (
    .A(_03066_),
    .B(_03153_),
    .C(_03064_),
    .Y(_03155_)
  );
  OAI22X1 _08609_ (
    .A(_02998_),
    .B(_03064_),
    .C(_03154_),
    .D(_03155_),
    .Y(_02032_)
  );
  AOI22X1 _08610_ (
    .A(execution_unit_0.register_file_0.r1_5_ ),
    .B(_03031_),
    .C(_03052_),
    .D(execution_unit_0.register_file_0.r15_5_ ),
    .Y(_03156_)
  );
  AOI22X1 _08611_ (
    .A(execution_unit_0.register_file_0.r9_5_ ),
    .B(_03025_),
    .C(_03027_),
    .D(execution_unit_0.register_file_0.r3_5_ ),
    .Y(_03157_)
  );
  NAND2X1 _08612_ (
    .A(_03156_),
    .B(_03157_),
    .Y(_03158_)
  );
  AOI22X1 _08613_ (
    .A(execution_unit_0.register_file_0.r10_5_ ),
    .B(_03044_),
    .C(_03047_),
    .D(execution_unit_0.register_file_0.r7_5_ ),
    .Y(_03159_)
  );
  AOI22X1 _08614_ (
    .A(execution_unit_0.register_file_0.r13_5_ ),
    .B(_03038_),
    .C(_03054_),
    .D(execution_unit_0.register_file_0.r5_5_ ),
    .Y(_03160_)
  );
  NAND2X1 _08615_ (
    .A(_03159_),
    .B(_03160_),
    .Y(_03161_)
  );
  NOR2X1 _08616_ (
    .A(_03158_),
    .B(_03161_),
    .Y(_03162_)
  );
  AOI22X1 _08617_ (
    .A(execution_unit_0.register_file_0.r8_5_ ),
    .B(_03034_),
    .C(_03049_),
    .D(dbg_0.UNUSED_pc_5_ ),
    .Y(_03163_)
  );
  AOI22X1 _08618_ (
    .A(execution_unit_0.register_file_0.r11_5_ ),
    .B(_03023_),
    .C(_03029_),
    .D(execution_unit_0.register_file_0.r12_5_ ),
    .Y(_03164_)
  );
  NAND2X1 _08619_ (
    .A(_03163_),
    .B(_03164_),
    .Y(_03165_)
  );
  AOI22X1 _08620_ (
    .A(execution_unit_0.register_file_0.r6_5_ ),
    .B(_03021_),
    .C(_03041_),
    .D(execution_unit_0.register_file_0.r4_5_ ),
    .Y(_03166_)
  );
  AOI22X1 _08621_ (
    .A(clock_module_0.oscoff ),
    .B(_03033_),
    .C(_03036_),
    .D(execution_unit_0.register_file_0.r14_5_ ),
    .Y(_03167_)
  );
  NAND2X1 _08622_ (
    .A(_03166_),
    .B(_03167_),
    .Y(_03168_)
  );
  NOR2X1 _08623_ (
    .A(_03165_),
    .B(_03168_),
    .Y(_03169_)
  );
  NAND2X1 _08624_ (
    .A(_03162_),
    .B(_03169_),
    .Y(execution_unit_0.reg_src_5_ )
  );
  NAND3X1 _08625_ (
    .A(_03133_),
    .B(execution_unit_0.reg_src_4_ ),
    .C(execution_unit_0.reg_src_5_ ),
    .Y(_03170_)
  );
  XNOR2X1 _08626_ (
    .A(_03152_),
    .B(execution_unit_0.reg_src_5_ ),
    .Y(_03171_)
  );
  NOR2X1 _08627_ (
    .A(execution_unit_0.register_file_0.r14_5_ ),
    .B(_03065_),
    .Y(_03172_)
  );
  OAI21X1 _08628_ (
    .A(_03066_),
    .B(_03171_),
    .C(_03064_),
    .Y(_03173_)
  );
  OAI22X1 _08629_ (
    .A(_03000_),
    .B(_03064_),
    .C(_03172_),
    .D(_03173_),
    .Y(_02033_)
  );
  AOI22X1 _08630_ (
    .A(execution_unit_0.register_file_0.r6_6_ ),
    .B(_03021_),
    .C(_03047_),
    .D(execution_unit_0.register_file_0.r7_6_ ),
    .Y(_03174_)
  );
  AOI22X1 _08631_ (
    .A(execution_unit_0.register_file_0.r1_6_ ),
    .B(_03031_),
    .C(_03036_),
    .D(execution_unit_0.register_file_0.r14_6_ ),
    .Y(_03175_)
  );
  AND2X1 _08632_ (
    .A(_03174_),
    .B(_03175_),
    .Y(_03176_)
  );
  AOI22X1 _08633_ (
    .A(execution_unit_0.register_file_0.r11_6_ ),
    .B(_03023_),
    .C(_03038_),
    .D(execution_unit_0.register_file_0.r13_6_ ),
    .Y(_03177_)
  );
  AOI22X1 _08634_ (
    .A(execution_unit_0.register_file_0.r3_6_ ),
    .B(_03027_),
    .C(_03054_),
    .D(execution_unit_0.register_file_0.r5_6_ ),
    .Y(_03178_)
  );
  NAND3X1 _08635_ (
    .A(_03176_),
    .B(_03177_),
    .C(_03178_),
    .Y(_03179_)
  );
  AOI22X1 _08636_ (
    .A(execution_unit_0.register_file_0.r4_6_ ),
    .B(_03041_),
    .C(_03052_),
    .D(execution_unit_0.register_file_0.r15_6_ ),
    .Y(_03180_)
  );
  INVX1 _08637_ (
    .A(_03180_),
    .Y(_03181_)
  );
  AOI21X1 _08638_ (
    .A(execution_unit_0.register_file_0.r9_6_ ),
    .B(_03025_),
    .C(_03181_),
    .Y(_03182_)
  );
  AOI22X1 _08639_ (
    .A(execution_unit_0.register_file_0.r10_6_ ),
    .B(_03044_),
    .C(_03049_),
    .D(dbg_0.UNUSED_pc_6_ ),
    .Y(_03183_)
  );
  AOI22X1 _08640_ (
    .A(execution_unit_0.register_file_0.r12_6_ ),
    .B(_03029_),
    .C(_03034_),
    .D(execution_unit_0.register_file_0.r8_6_ ),
    .Y(_03184_)
  );
  NAND3X1 _08641_ (
    .A(_03182_),
    .B(_03183_),
    .C(_03184_),
    .Y(_03185_)
  );
  NOR2X1 _08642_ (
    .A(_03179_),
    .B(_03185_),
    .Y(_03186_)
  );
  INVX1 _08643_ (
    .A(_03186_),
    .Y(execution_unit_0.reg_src_6_ )
  );
  NOR2X1 _08644_ (
    .A(_03170_),
    .B(_03186_),
    .Y(_03187_)
  );
  XNOR2X1 _08645_ (
    .A(_03170_),
    .B(execution_unit_0.reg_src_6_ ),
    .Y(_03188_)
  );
  NOR2X1 _08646_ (
    .A(execution_unit_0.register_file_0.r14_6_ ),
    .B(_03065_),
    .Y(_03189_)
  );
  OAI21X1 _08647_ (
    .A(_03066_),
    .B(_03188_),
    .C(_03064_),
    .Y(_03190_)
  );
  OAI22X1 _08648_ (
    .A(_03002_),
    .B(_03064_),
    .C(_03189_),
    .D(_03190_),
    .Y(_02034_)
  );
  AOI22X1 _08649_ (
    .A(execution_unit_0.register_file_0.r9_7_ ),
    .B(_03025_),
    .C(_03049_),
    .D(dbg_0.UNUSED_pc_7_ ),
    .Y(_03191_)
  );
  AOI22X1 _08650_ (
    .A(execution_unit_0.register_file_0.r7_7_ ),
    .B(_03047_),
    .C(_03054_),
    .D(execution_unit_0.register_file_0.r5_7_ ),
    .Y(_03192_)
  );
  NAND2X1 _08651_ (
    .A(_03191_),
    .B(_03192_),
    .Y(_03193_)
  );
  AOI22X1 _08652_ (
    .A(execution_unit_0.register_file_0.r1_7_ ),
    .B(_03031_),
    .C(_03038_),
    .D(execution_unit_0.register_file_0.r13_7_ ),
    .Y(_03194_)
  );
  AOI22X1 _08653_ (
    .A(execution_unit_0.register_file_0.r8_7_ ),
    .B(_03034_),
    .C(_03052_),
    .D(execution_unit_0.register_file_0.r15_7_ ),
    .Y(_03195_)
  );
  NAND2X1 _08654_ (
    .A(_03194_),
    .B(_03195_),
    .Y(_03196_)
  );
  NOR2X1 _08655_ (
    .A(_03193_),
    .B(_03196_),
    .Y(_03197_)
  );
  AOI22X1 _08656_ (
    .A(execution_unit_0.register_file_0.r6_7_ ),
    .B(_03021_),
    .C(_03023_),
    .D(execution_unit_0.register_file_0.r11_7_ ),
    .Y(_03198_)
  );
  AOI22X1 _08657_ (
    .A(execution_unit_0.register_file_0.r12_7_ ),
    .B(_03029_),
    .C(_03044_),
    .D(execution_unit_0.register_file_0.r10_7_ ),
    .Y(_03199_)
  );
  NAND2X1 _08658_ (
    .A(_03198_),
    .B(_03199_),
    .Y(_03200_)
  );
  AOI22X1 _08659_ (
    .A(execution_unit_0.register_file_0.r3_7_ ),
    .B(_03027_),
    .C(_03036_),
    .D(execution_unit_0.register_file_0.r14_7_ ),
    .Y(_03201_)
  );
  AOI22X1 _08660_ (
    .A(clock_module_0.scg1 ),
    .B(_03033_),
    .C(_03041_),
    .D(execution_unit_0.register_file_0.r4_7_ ),
    .Y(_03202_)
  );
  NAND2X1 _08661_ (
    .A(_03201_),
    .B(_03202_),
    .Y(_03203_)
  );
  NOR2X1 _08662_ (
    .A(_03200_),
    .B(_03203_),
    .Y(_03204_)
  );
  NAND2X1 _08663_ (
    .A(_03197_),
    .B(_03204_),
    .Y(execution_unit_0.reg_src_7_ )
  );
  INVX1 _08664_ (
    .A(execution_unit_0.reg_src_7_ ),
    .Y(_03205_)
  );
  NOR3X1 _08665_ (
    .A(_03170_),
    .B(_03186_),
    .C(_03205_),
    .Y(_03206_)
  );
  NOR2X1 _08666_ (
    .A(_03187_),
    .B(execution_unit_0.reg_src_7_ ),
    .Y(_03207_)
  );
  NOR2X1 _08667_ (
    .A(_03206_),
    .B(_03207_),
    .Y(_03208_)
  );
  NOR2X1 _08668_ (
    .A(execution_unit_0.register_file_0.r14_7_ ),
    .B(_03065_),
    .Y(_03209_)
  );
  OAI21X1 _08669_ (
    .A(_03066_),
    .B(_03208_),
    .C(_03064_),
    .Y(_03210_)
  );
  OAI22X1 _08670_ (
    .A(_03004_),
    .B(_03064_),
    .C(_03209_),
    .D(_03210_),
    .Y(_02035_)
  );
  NAND2X1 _08671_ (
    .A(_02982_),
    .B(execution_unit_0.alu_0.alu_out_8_ ),
    .Y(_03211_)
  );
  INVX1 _08672_ (
    .A(_03211_),
    .Y(execution_unit_0.pc_sw_8_ )
  );
  AOI22X1 _08673_ (
    .A(execution_unit_0.register_file_0.r11_8_ ),
    .B(_03023_),
    .C(_03034_),
    .D(execution_unit_0.register_file_0.r8_8_ ),
    .Y(_03212_)
  );
  AOI22X1 _08674_ (
    .A(execution_unit_0.register_file_0.r1_8_ ),
    .B(_03031_),
    .C(_03033_),
    .D(execution_unit_0.alu_0.status_3_ ),
    .Y(_03213_)
  );
  NAND2X1 _08675_ (
    .A(_03212_),
    .B(_03213_),
    .Y(_03214_)
  );
  AOI22X1 _08676_ (
    .A(dbg_0.UNUSED_pc_8_ ),
    .B(_03049_),
    .C(_03052_),
    .D(execution_unit_0.register_file_0.r15_8_ ),
    .Y(_03215_)
  );
  AOI22X1 _08677_ (
    .A(execution_unit_0.register_file_0.r14_8_ ),
    .B(_03036_),
    .C(_03047_),
    .D(execution_unit_0.register_file_0.r7_8_ ),
    .Y(_03216_)
  );
  NAND2X1 _08678_ (
    .A(_03215_),
    .B(_03216_),
    .Y(_03217_)
  );
  NOR2X1 _08679_ (
    .A(_03214_),
    .B(_03217_),
    .Y(_03218_)
  );
  AOI22X1 _08680_ (
    .A(execution_unit_0.register_file_0.r6_8_ ),
    .B(_03021_),
    .C(_03041_),
    .D(execution_unit_0.register_file_0.r4_8_ ),
    .Y(_03219_)
  );
  AOI22X1 _08681_ (
    .A(execution_unit_0.register_file_0.r13_8_ ),
    .B(_03038_),
    .C(_03054_),
    .D(execution_unit_0.register_file_0.r5_8_ ),
    .Y(_03220_)
  );
  NAND2X1 _08682_ (
    .A(_03219_),
    .B(_03220_),
    .Y(_03221_)
  );
  AOI22X1 _08683_ (
    .A(execution_unit_0.register_file_0.r3_8_ ),
    .B(_03027_),
    .C(_03029_),
    .D(execution_unit_0.register_file_0.r12_8_ ),
    .Y(_03222_)
  );
  AOI22X1 _08684_ (
    .A(execution_unit_0.register_file_0.r9_8_ ),
    .B(_03025_),
    .C(_03044_),
    .D(execution_unit_0.register_file_0.r10_8_ ),
    .Y(_03223_)
  );
  NAND2X1 _08685_ (
    .A(_03222_),
    .B(_03223_),
    .Y(_03224_)
  );
  NOR2X1 _08686_ (
    .A(_03221_),
    .B(_03224_),
    .Y(_03225_)
  );
  NAND2X1 _08687_ (
    .A(_03218_),
    .B(_03225_),
    .Y(execution_unit_0.reg_src_8_ )
  );
  NAND2X1 _08688_ (
    .A(_03206_),
    .B(execution_unit_0.reg_src_8_ ),
    .Y(_03226_)
  );
  XOR2X1 _08689_ (
    .A(_03206_),
    .B(execution_unit_0.reg_src_8_ ),
    .Y(_03227_)
  );
  OAI21X1 _08690_ (
    .A(_03066_),
    .B(_03227_),
    .C(_03064_),
    .Y(_03228_)
  );
  INVX1 _08691_ (
    .A(_03228_),
    .Y(_03229_)
  );
  OAI21X1 _08692_ (
    .A(execution_unit_0.register_file_0.r14_8_ ),
    .B(_03065_),
    .C(_03229_),
    .Y(_03230_)
  );
  OAI21X1 _08693_ (
    .A(_03064_),
    .B(_03211_),
    .C(_03230_),
    .Y(_02036_)
  );
  NAND2X1 _08694_ (
    .A(_02982_),
    .B(execution_unit_0.alu_0.alu_out_9_ ),
    .Y(_03231_)
  );
  INVX1 _08695_ (
    .A(_03231_),
    .Y(execution_unit_0.pc_sw_9_ )
  );
  AOI22X1 _08696_ (
    .A(execution_unit_0.register_file_0.r3_9_ ),
    .B(_03027_),
    .C(_03029_),
    .D(execution_unit_0.register_file_0.r12_9_ ),
    .Y(_03232_)
  );
  OAI21X1 _08697_ (
    .A(_03007_),
    .B(_03039_),
    .C(_03232_),
    .Y(_03233_)
  );
  AOI21X1 _08698_ (
    .A(execution_unit_0.register_file_0.r5_9_ ),
    .B(_03054_),
    .C(_03233_),
    .Y(_03234_)
  );
  AOI22X1 _08699_ (
    .A(execution_unit_0.register_file_0.r11_9_ ),
    .B(_03023_),
    .C(_03047_),
    .D(execution_unit_0.register_file_0.r7_9_ ),
    .Y(_03235_)
  );
  AOI22X1 _08700_ (
    .A(execution_unit_0.register_file_0.r9_9_ ),
    .B(_03025_),
    .C(_03049_),
    .D(dbg_0.UNUSED_pc_9_ ),
    .Y(_03236_)
  );
  AND2X1 _08701_ (
    .A(_03235_),
    .B(_03236_),
    .Y(_03237_)
  );
  AOI22X1 _08702_ (
    .A(execution_unit_0.register_file_0.r1_9_ ),
    .B(_03031_),
    .C(_03052_),
    .D(execution_unit_0.register_file_0.r15_9_ ),
    .Y(_03238_)
  );
  AOI22X1 _08703_ (
    .A(execution_unit_0.register_file_0.r4_9_ ),
    .B(_03041_),
    .C(_03044_),
    .D(execution_unit_0.register_file_0.r10_9_ ),
    .Y(_03239_)
  );
  AOI22X1 _08704_ (
    .A(execution_unit_0.register_file_0.r8_9_ ),
    .B(_03034_),
    .C(_03036_),
    .D(execution_unit_0.register_file_0.r14_9_ ),
    .Y(_03240_)
  );
  NAND3X1 _08705_ (
    .A(_03238_),
    .B(_03239_),
    .C(_03240_),
    .Y(_03241_)
  );
  AOI21X1 _08706_ (
    .A(execution_unit_0.register_file_0.r6_9_ ),
    .B(_03021_),
    .C(_03241_),
    .Y(_03242_)
  );
  NAND3X1 _08707_ (
    .A(_03234_),
    .B(_03237_),
    .C(_03242_),
    .Y(execution_unit_0.reg_src_9_ )
  );
  NAND3X1 _08708_ (
    .A(_03206_),
    .B(execution_unit_0.reg_src_8_ ),
    .C(execution_unit_0.reg_src_9_ ),
    .Y(_03243_)
  );
  XNOR2X1 _08709_ (
    .A(_03226_),
    .B(execution_unit_0.reg_src_9_ ),
    .Y(_03244_)
  );
  OAI21X1 _08710_ (
    .A(_03066_),
    .B(_03244_),
    .C(_03064_),
    .Y(_03245_)
  );
  INVX1 _08711_ (
    .A(_03245_),
    .Y(_03246_)
  );
  OAI21X1 _08712_ (
    .A(execution_unit_0.register_file_0.r14_9_ ),
    .B(_03065_),
    .C(_03246_),
    .Y(_03247_)
  );
  OAI21X1 _08713_ (
    .A(_03064_),
    .B(_03231_),
    .C(_03247_),
    .Y(_02037_)
  );
  NAND2X1 _08714_ (
    .A(_02982_),
    .B(execution_unit_0.alu_0.alu_out_10_ ),
    .Y(_03248_)
  );
  INVX1 _08715_ (
    .A(_03248_),
    .Y(execution_unit_0.pc_sw_10_ )
  );
  NAND2X1 _08716_ (
    .A(execution_unit_0.register_file_0.r6_10_ ),
    .B(_03021_),
    .Y(_03249_)
  );
  AOI22X1 _08717_ (
    .A(execution_unit_0.register_file_0.r13_10_ ),
    .B(_03038_),
    .C(_03054_),
    .D(execution_unit_0.register_file_0.r5_10_ ),
    .Y(_03250_)
  );
  OAI21X1 _08718_ (
    .A(_03008_),
    .B(_03042_),
    .C(_03250_),
    .Y(_03251_)
  );
  AOI22X1 _08719_ (
    .A(execution_unit_0.register_file_0.r3_10_ ),
    .B(_03027_),
    .C(_03044_),
    .D(execution_unit_0.register_file_0.r10_10_ ),
    .Y(_03252_)
  );
  AOI22X1 _08720_ (
    .A(execution_unit_0.register_file_0.r1_10_ ),
    .B(_03031_),
    .C(_03036_),
    .D(execution_unit_0.register_file_0.r14_10_ ),
    .Y(_03253_)
  );
  AOI22X1 _08721_ (
    .A(dbg_0.UNUSED_pc_10_ ),
    .B(_03049_),
    .C(_03052_),
    .D(execution_unit_0.register_file_0.r15_10_ ),
    .Y(_03254_)
  );
  NAND3X1 _08722_ (
    .A(_03252_),
    .B(_03253_),
    .C(_03254_),
    .Y(_03255_)
  );
  AOI21X1 _08723_ (
    .A(execution_unit_0.register_file_0.r8_10_ ),
    .B(_03034_),
    .C(_03255_),
    .Y(_03256_)
  );
  INVX1 _08724_ (
    .A(_03256_),
    .Y(_03257_)
  );
  AOI22X1 _08725_ (
    .A(execution_unit_0.register_file_0.r12_10_ ),
    .B(_03029_),
    .C(_03047_),
    .D(execution_unit_0.register_file_0.r7_10_ ),
    .Y(_03258_)
  );
  AOI22X1 _08726_ (
    .A(execution_unit_0.register_file_0.r11_10_ ),
    .B(_03023_),
    .C(_03025_),
    .D(execution_unit_0.register_file_0.r9_10_ ),
    .Y(_03259_)
  );
  NAND2X1 _08727_ (
    .A(_03249_),
    .B(_03259_),
    .Y(_03260_)
  );
  NOR2X1 _08728_ (
    .A(_03251_),
    .B(_03260_),
    .Y(_03261_)
  );
  NAND2X1 _08729_ (
    .A(_03258_),
    .B(_03261_),
    .Y(_03262_)
  );
  NOR2X1 _08730_ (
    .A(_03257_),
    .B(_03262_),
    .Y(_03263_)
  );
  INVX1 _08731_ (
    .A(_03263_),
    .Y(execution_unit_0.reg_src_10_ )
  );
  NOR2X1 _08732_ (
    .A(_03243_),
    .B(_03263_),
    .Y(_03264_)
  );
  XNOR2X1 _08733_ (
    .A(_03243_),
    .B(_03263_),
    .Y(_03265_)
  );
  AOI21X1 _08734_ (
    .A(_03065_),
    .B(_03265_),
    .C(_03063_),
    .Y(_03266_)
  );
  OAI21X1 _08735_ (
    .A(execution_unit_0.register_file_0.r14_10_ ),
    .B(_03065_),
    .C(_03266_),
    .Y(_03267_)
  );
  OAI21X1 _08736_ (
    .A(_03064_),
    .B(_03248_),
    .C(_03267_),
    .Y(_02023_)
  );
  NAND2X1 _08737_ (
    .A(_02982_),
    .B(execution_unit_0.alu_0.alu_out_11_ ),
    .Y(_03268_)
  );
  INVX1 _08738_ (
    .A(_03268_),
    .Y(execution_unit_0.pc_sw_11_ )
  );
  NAND2X1 _08739_ (
    .A(execution_unit_0.register_file_0.r4_11_ ),
    .B(_03041_),
    .Y(_03269_)
  );
  NAND2X1 _08740_ (
    .A(execution_unit_0.register_file_0.r10_11_ ),
    .B(_03044_),
    .Y(_03270_)
  );
  AOI22X1 _08741_ (
    .A(execution_unit_0.register_file_0.r9_11_ ),
    .B(_03025_),
    .C(_03038_),
    .D(execution_unit_0.register_file_0.r13_11_ ),
    .Y(_03271_)
  );
  AOI22X1 _08742_ (
    .A(execution_unit_0.register_file_0.r14_11_ ),
    .B(_03036_),
    .C(_03052_),
    .D(execution_unit_0.register_file_0.r15_11_ ),
    .Y(_03272_)
  );
  AOI22X1 _08743_ (
    .A(execution_unit_0.register_file_0.r6_11_ ),
    .B(_03021_),
    .C(_03029_),
    .D(execution_unit_0.register_file_0.r12_11_ ),
    .Y(_03273_)
  );
  NAND2X1 _08744_ (
    .A(_03272_),
    .B(_03273_),
    .Y(_03274_)
  );
  AOI21X1 _08745_ (
    .A(execution_unit_0.register_file_0.r8_11_ ),
    .B(_03034_),
    .C(_03274_),
    .Y(_03275_)
  );
  NAND3X1 _08746_ (
    .A(_03269_),
    .B(_03270_),
    .C(_03271_),
    .Y(_03276_)
  );
  AOI22X1 _08747_ (
    .A(execution_unit_0.register_file_0.r7_11_ ),
    .B(_03047_),
    .C(_03054_),
    .D(execution_unit_0.register_file_0.r5_11_ ),
    .Y(_03277_)
  );
  AOI22X1 _08748_ (
    .A(execution_unit_0.register_file_0.r11_11_ ),
    .B(_03023_),
    .C(_03027_),
    .D(execution_unit_0.register_file_0.r3_11_ ),
    .Y(_03278_)
  );
  AOI22X1 _08749_ (
    .A(execution_unit_0.register_file_0.r1_11_ ),
    .B(_03031_),
    .C(_03049_),
    .D(dbg_0.UNUSED_pc_11_ ),
    .Y(_03279_)
  );
  NAND3X1 _08750_ (
    .A(_03277_),
    .B(_03278_),
    .C(_03279_),
    .Y(_03280_)
  );
  NOR2X1 _08751_ (
    .A(_03276_),
    .B(_03280_),
    .Y(_03281_)
  );
  NAND2X1 _08752_ (
    .A(_03275_),
    .B(_03281_),
    .Y(execution_unit_0.reg_src_11_ )
  );
  INVX1 _08753_ (
    .A(execution_unit_0.reg_src_11_ ),
    .Y(_03282_)
  );
  NOR3X1 _08754_ (
    .A(_03243_),
    .B(_03263_),
    .C(_03282_),
    .Y(_03283_)
  );
  XNOR2X1 _08755_ (
    .A(_03264_),
    .B(_03282_),
    .Y(_03284_)
  );
  OAI21X1 _08756_ (
    .A(_03066_),
    .B(_03284_),
    .C(_03064_),
    .Y(_03285_)
  );
  INVX1 _08757_ (
    .A(_03285_),
    .Y(_03286_)
  );
  OAI21X1 _08758_ (
    .A(execution_unit_0.register_file_0.r14_11_ ),
    .B(_03065_),
    .C(_03286_),
    .Y(_03287_)
  );
  OAI21X1 _08759_ (
    .A(_03064_),
    .B(_03268_),
    .C(_03287_),
    .Y(_02024_)
  );
  NAND2X1 _08760_ (
    .A(_02982_),
    .B(execution_unit_0.alu_0.alu_out_12_ ),
    .Y(_03288_)
  );
  INVX1 _08761_ (
    .A(_03288_),
    .Y(execution_unit_0.pc_sw_12_ )
  );
  AOI22X1 _08762_ (
    .A(execution_unit_0.register_file_0.r13_12_ ),
    .B(_03038_),
    .C(_03044_),
    .D(execution_unit_0.register_file_0.r10_12_ ),
    .Y(_03289_)
  );
  AOI22X1 _08763_ (
    .A(execution_unit_0.register_file_0.r6_12_ ),
    .B(_03021_),
    .C(_03027_),
    .D(execution_unit_0.register_file_0.r3_12_ ),
    .Y(_03290_)
  );
  AND2X1 _08764_ (
    .A(_03289_),
    .B(_03290_),
    .Y(_03291_)
  );
  AOI22X1 _08765_ (
    .A(execution_unit_0.register_file_0.r8_12_ ),
    .B(_03034_),
    .C(_03036_),
    .D(execution_unit_0.register_file_0.r14_12_ ),
    .Y(_03292_)
  );
  AOI22X1 _08766_ (
    .A(execution_unit_0.register_file_0.r1_12_ ),
    .B(_03031_),
    .C(_03049_),
    .D(dbg_0.UNUSED_pc_12_ ),
    .Y(_03293_)
  );
  NAND3X1 _08767_ (
    .A(_03291_),
    .B(_03292_),
    .C(_03293_),
    .Y(_03294_)
  );
  AOI22X1 _08768_ (
    .A(execution_unit_0.register_file_0.r15_12_ ),
    .B(_03052_),
    .C(_03054_),
    .D(execution_unit_0.register_file_0.r5_12_ ),
    .Y(_03295_)
  );
  INVX1 _08769_ (
    .A(_03295_),
    .Y(_03296_)
  );
  AOI21X1 _08770_ (
    .A(execution_unit_0.register_file_0.r11_12_ ),
    .B(_03023_),
    .C(_03296_),
    .Y(_03297_)
  );
  AOI22X1 _08771_ (
    .A(execution_unit_0.register_file_0.r9_12_ ),
    .B(_03025_),
    .C(_03041_),
    .D(execution_unit_0.register_file_0.r4_12_ ),
    .Y(_03298_)
  );
  AOI22X1 _08772_ (
    .A(execution_unit_0.register_file_0.r12_12_ ),
    .B(_03029_),
    .C(_03047_),
    .D(execution_unit_0.register_file_0.r7_12_ ),
    .Y(_03299_)
  );
  NAND3X1 _08773_ (
    .A(_03297_),
    .B(_03298_),
    .C(_03299_),
    .Y(_03300_)
  );
  OR2X1 _08774_ (
    .A(_03294_),
    .B(_03300_),
    .Y(execution_unit_0.reg_src_12_ )
  );
  OAI21X1 _08775_ (
    .A(_03294_),
    .B(_03300_),
    .C(_03283_),
    .Y(_03301_)
  );
  XOR2X1 _08776_ (
    .A(_03283_),
    .B(execution_unit_0.reg_src_12_ ),
    .Y(_03302_)
  );
  OAI21X1 _08777_ (
    .A(execution_unit_0.register_file_0.r14_12_ ),
    .B(_03065_),
    .C(_03064_),
    .Y(_03303_)
  );
  INVX1 _08778_ (
    .A(_03303_),
    .Y(_03304_)
  );
  OAI21X1 _08779_ (
    .A(_03066_),
    .B(_03302_),
    .C(_03304_),
    .Y(_03305_)
  );
  OAI21X1 _08780_ (
    .A(_03064_),
    .B(_03288_),
    .C(_03305_),
    .Y(_02025_)
  );
  NAND2X1 _08781_ (
    .A(_02982_),
    .B(execution_unit_0.alu_0.alu_out_13_ ),
    .Y(_03306_)
  );
  INVX1 _08782_ (
    .A(_03306_),
    .Y(execution_unit_0.pc_sw_13_ )
  );
  NAND2X1 _08783_ (
    .A(execution_unit_0.register_file_0.r13_13_ ),
    .B(_03038_),
    .Y(_03307_)
  );
  NAND2X1 _08784_ (
    .A(dbg_0.UNUSED_pc_13_ ),
    .B(_03049_),
    .Y(_03308_)
  );
  AOI22X1 _08785_ (
    .A(execution_unit_0.register_file_0.r6_13_ ),
    .B(_03021_),
    .C(_03052_),
    .D(execution_unit_0.register_file_0.r15_13_ ),
    .Y(_03309_)
  );
  AOI22X1 _08786_ (
    .A(execution_unit_0.register_file_0.r8_13_ ),
    .B(_03034_),
    .C(_03044_),
    .D(execution_unit_0.register_file_0.r10_13_ ),
    .Y(_03310_)
  );
  AOI22X1 _08787_ (
    .A(execution_unit_0.register_file_0.r12_13_ ),
    .B(_03029_),
    .C(_03036_),
    .D(execution_unit_0.register_file_0.r14_13_ ),
    .Y(_03311_)
  );
  AOI22X1 _08788_ (
    .A(execution_unit_0.register_file_0.r7_13_ ),
    .B(_03047_),
    .C(_03054_),
    .D(execution_unit_0.register_file_0.r5_13_ ),
    .Y(_03312_)
  );
  AOI22X1 _08789_ (
    .A(execution_unit_0.register_file_0.r9_13_ ),
    .B(_03025_),
    .C(_03031_),
    .D(execution_unit_0.register_file_0.r1_13_ ),
    .Y(_03313_)
  );
  NAND2X1 _08790_ (
    .A(_03312_),
    .B(_03313_),
    .Y(_03314_)
  );
  AOI21X1 _08791_ (
    .A(execution_unit_0.register_file_0.r11_13_ ),
    .B(_03023_),
    .C(_03314_),
    .Y(_03315_)
  );
  NAND3X1 _08792_ (
    .A(_03307_),
    .B(_03308_),
    .C(_03311_),
    .Y(_03316_)
  );
  AOI22X1 _08793_ (
    .A(execution_unit_0.register_file_0.r3_13_ ),
    .B(_03027_),
    .C(_03041_),
    .D(execution_unit_0.register_file_0.r4_13_ ),
    .Y(_03317_)
  );
  NAND3X1 _08794_ (
    .A(_03309_),
    .B(_03310_),
    .C(_03317_),
    .Y(_03318_)
  );
  NOR2X1 _08795_ (
    .A(_03316_),
    .B(_03318_),
    .Y(_03319_)
  );
  NAND2X1 _08796_ (
    .A(_03315_),
    .B(_03319_),
    .Y(execution_unit_0.reg_src_13_ )
  );
  NAND3X1 _08797_ (
    .A(_03283_),
    .B(execution_unit_0.reg_src_12_ ),
    .C(execution_unit_0.reg_src_13_ ),
    .Y(_03320_)
  );
  XNOR2X1 _08798_ (
    .A(_03301_),
    .B(execution_unit_0.reg_src_13_ ),
    .Y(_03321_)
  );
  OAI21X1 _08799_ (
    .A(execution_unit_0.register_file_0.r14_13_ ),
    .B(_03065_),
    .C(_03064_),
    .Y(_03322_)
  );
  INVX1 _08800_ (
    .A(_03322_),
    .Y(_03323_)
  );
  OAI21X1 _08801_ (
    .A(_03066_),
    .B(_03321_),
    .C(_03323_),
    .Y(_03324_)
  );
  OAI21X1 _08802_ (
    .A(_03064_),
    .B(_03306_),
    .C(_03324_),
    .Y(_02026_)
  );
  NAND2X1 _08803_ (
    .A(_02982_),
    .B(execution_unit_0.alu_0.alu_out_14_ ),
    .Y(_03325_)
  );
  INVX1 _08804_ (
    .A(_03325_),
    .Y(execution_unit_0.pc_sw_14_ )
  );
  NAND2X1 _08805_ (
    .A(execution_unit_0.register_file_0.r14_14_ ),
    .B(_03036_),
    .Y(_03326_)
  );
  AOI22X1 _08806_ (
    .A(execution_unit_0.register_file_0.r13_14_ ),
    .B(_03038_),
    .C(_03052_),
    .D(execution_unit_0.register_file_0.r15_14_ ),
    .Y(_03327_)
  );
  NAND2X1 _08807_ (
    .A(_03326_),
    .B(_03327_),
    .Y(_03328_)
  );
  AOI22X1 _08808_ (
    .A(execution_unit_0.register_file_0.r8_14_ ),
    .B(_03034_),
    .C(_03047_),
    .D(execution_unit_0.register_file_0.r7_14_ ),
    .Y(_03329_)
  );
  AOI22X1 _08809_ (
    .A(execution_unit_0.register_file_0.r6_14_ ),
    .B(_03021_),
    .C(_03049_),
    .D(dbg_0.UNUSED_pc_14_ ),
    .Y(_03330_)
  );
  AOI22X1 _08810_ (
    .A(execution_unit_0.register_file_0.r4_14_ ),
    .B(_03041_),
    .C(_03054_),
    .D(execution_unit_0.register_file_0.r5_14_ ),
    .Y(_03331_)
  );
  NAND3X1 _08811_ (
    .A(_03329_),
    .B(_03330_),
    .C(_03331_),
    .Y(_03332_)
  );
  AOI21X1 _08812_ (
    .A(execution_unit_0.register_file_0.r9_14_ ),
    .B(_03025_),
    .C(_03332_),
    .Y(_03333_)
  );
  AOI22X1 _08813_ (
    .A(execution_unit_0.register_file_0.r3_14_ ),
    .B(_03027_),
    .C(_03031_),
    .D(execution_unit_0.register_file_0.r1_14_ ),
    .Y(_03334_)
  );
  AOI22X1 _08814_ (
    .A(execution_unit_0.register_file_0.r11_14_ ),
    .B(_03023_),
    .C(_03029_),
    .D(execution_unit_0.register_file_0.r12_14_ ),
    .Y(_03335_)
  );
  OAI21X1 _08815_ (
    .A(_03013_),
    .B(_03045_),
    .C(_03335_),
    .Y(_03336_)
  );
  NOR2X1 _08816_ (
    .A(_03328_),
    .B(_03336_),
    .Y(_03337_)
  );
  NAND3X1 _08817_ (
    .A(_03333_),
    .B(_03334_),
    .C(_03337_),
    .Y(execution_unit_0.reg_src_14_ )
  );
  INVX1 _08818_ (
    .A(execution_unit_0.reg_src_14_ ),
    .Y(_03338_)
  );
  NOR2X1 _08819_ (
    .A(_03320_),
    .B(_03338_),
    .Y(_03339_)
  );
  XNOR2X1 _08820_ (
    .A(_03320_),
    .B(execution_unit_0.reg_src_14_ ),
    .Y(_02191_)
  );
  OAI21X1 _08821_ (
    .A(execution_unit_0.register_file_0.r14_14_ ),
    .B(_03065_),
    .C(_03064_),
    .Y(_02192_)
  );
  INVX1 _08822_ (
    .A(_02192_),
    .Y(_02193_)
  );
  OAI21X1 _08823_ (
    .A(_03066_),
    .B(_02191_),
    .C(_02193_),
    .Y(_02194_)
  );
  OAI21X1 _08824_ (
    .A(_03064_),
    .B(_03325_),
    .C(_02194_),
    .Y(_02027_)
  );
  NAND2X1 _08825_ (
    .A(_02982_),
    .B(execution_unit_0.alu_0.alu_out_15_ ),
    .Y(_02195_)
  );
  INVX1 _08826_ (
    .A(_02195_),
    .Y(execution_unit_0.pc_sw_15_ )
  );
  AOI22X1 _08827_ (
    .A(execution_unit_0.register_file_0.r3_15_ ),
    .B(_03027_),
    .C(_03052_),
    .D(execution_unit_0.register_file_0.r15_15_ ),
    .Y(_02196_)
  );
  NAND2X1 _08828_ (
    .A(execution_unit_0.register_file_0.r12_15_ ),
    .B(_03029_),
    .Y(_02197_)
  );
  OAI21X1 _08829_ (
    .A(_03014_),
    .B(_03039_),
    .C(_02196_),
    .Y(_02198_)
  );
  AOI21X1 _08830_ (
    .A(execution_unit_0.register_file_0.r8_15_ ),
    .B(_03034_),
    .C(_02198_),
    .Y(_02199_)
  );
  AOI22X1 _08831_ (
    .A(execution_unit_0.register_file_0.r1_15_ ),
    .B(_03031_),
    .C(_03049_),
    .D(dbg_0.UNUSED_pc_15_ ),
    .Y(_02200_)
  );
  AOI22X1 _08832_ (
    .A(execution_unit_0.register_file_0.r6_15_ ),
    .B(_03021_),
    .C(_03054_),
    .D(execution_unit_0.register_file_0.r5_15_ ),
    .Y(_02201_)
  );
  NAND2X1 _08833_ (
    .A(_02200_),
    .B(_02201_),
    .Y(_02202_)
  );
  AOI21X1 _08834_ (
    .A(execution_unit_0.register_file_0.r4_15_ ),
    .B(_03041_),
    .C(_02202_),
    .Y(_02203_)
  );
  AOI22X1 _08835_ (
    .A(execution_unit_0.register_file_0.r14_15_ ),
    .B(_03036_),
    .C(_03044_),
    .D(execution_unit_0.register_file_0.r10_15_ ),
    .Y(_02204_)
  );
  AOI22X1 _08836_ (
    .A(execution_unit_0.register_file_0.r9_15_ ),
    .B(_03025_),
    .C(_03047_),
    .D(execution_unit_0.register_file_0.r7_15_ ),
    .Y(_02205_)
  );
  NAND3X1 _08837_ (
    .A(_02197_),
    .B(_02204_),
    .C(_02205_),
    .Y(_02206_)
  );
  AOI21X1 _08838_ (
    .A(execution_unit_0.register_file_0.r11_15_ ),
    .B(_03023_),
    .C(_02206_),
    .Y(_02207_)
  );
  NAND3X1 _08839_ (
    .A(_02199_),
    .B(_02203_),
    .C(_02207_),
    .Y(execution_unit_0.reg_src_15_ )
  );
  XOR2X1 _08840_ (
    .A(_03339_),
    .B(execution_unit_0.reg_src_15_ ),
    .Y(_02208_)
  );
  OAI21X1 _08841_ (
    .A(execution_unit_0.register_file_0.r14_15_ ),
    .B(_03065_),
    .C(_03064_),
    .Y(_02209_)
  );
  INVX1 _08842_ (
    .A(_02209_),
    .Y(_02210_)
  );
  OAI21X1 _08843_ (
    .A(_03066_),
    .B(_02208_),
    .C(_02210_),
    .Y(_02211_)
  );
  OAI21X1 _08844_ (
    .A(_03064_),
    .B(_02195_),
    .C(_02211_),
    .Y(_02028_)
  );
  AND2X1 _08845_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_15_ ),
    .Y(_02212_)
  );
  NAND2X1 _08846_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_15_ ),
    .Y(_02213_)
  );
  AND2X1 _08847_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03052_),
    .Y(_02214_)
  );
  NAND2X1 _08848_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03052_),
    .Y(_02215_)
  );
  AOI21X1 _08849_ (
    .A(_03069_),
    .B(_02214_),
    .C(_02212_),
    .Y(_02216_)
  );
  OAI21X1 _08850_ (
    .A(execution_unit_0.register_file_0.r15_0_ ),
    .B(_02214_),
    .C(_02216_),
    .Y(_02217_)
  );
  OAI21X1 _08851_ (
    .A(_02984_),
    .B(_02213_),
    .C(_02217_),
    .Y(_02038_)
  );
  NOR2X1 _08852_ (
    .A(execution_unit_0.register_file_0.r15_1_ ),
    .B(_02214_),
    .Y(_02218_)
  );
  OAI21X1 _08853_ (
    .A(_03093_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02219_)
  );
  OAI22X1 _08854_ (
    .A(_02989_),
    .B(_02213_),
    .C(_02218_),
    .D(_02219_),
    .Y(_02045_)
  );
  AOI21X1 _08855_ (
    .A(_03112_),
    .B(_02214_),
    .C(_02212_),
    .Y(_02220_)
  );
  OAI21X1 _08856_ (
    .A(execution_unit_0.register_file_0.r15_2_ ),
    .B(_02214_),
    .C(_02220_),
    .Y(_02221_)
  );
  OAI21X1 _08857_ (
    .A(_02991_),
    .B(_02213_),
    .C(_02221_),
    .Y(_02046_)
  );
  NOR2X1 _08858_ (
    .A(execution_unit_0.register_file_0.r15_3_ ),
    .B(_02214_),
    .Y(_02222_)
  );
  OAI21X1 _08859_ (
    .A(_03135_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02223_)
  );
  OAI22X1 _08860_ (
    .A(_02995_),
    .B(_02213_),
    .C(_02222_),
    .D(_02223_),
    .Y(_02047_)
  );
  NOR2X1 _08861_ (
    .A(execution_unit_0.register_file_0.r15_4_ ),
    .B(_02214_),
    .Y(_02224_)
  );
  OAI21X1 _08862_ (
    .A(_03153_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02225_)
  );
  OAI22X1 _08863_ (
    .A(_02998_),
    .B(_02213_),
    .C(_02224_),
    .D(_02225_),
    .Y(_02048_)
  );
  NOR2X1 _08864_ (
    .A(execution_unit_0.register_file_0.r15_5_ ),
    .B(_02214_),
    .Y(_02226_)
  );
  OAI21X1 _08865_ (
    .A(_03171_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02227_)
  );
  OAI22X1 _08866_ (
    .A(_03000_),
    .B(_02213_),
    .C(_02226_),
    .D(_02227_),
    .Y(_02049_)
  );
  NOR2X1 _08867_ (
    .A(execution_unit_0.register_file_0.r15_6_ ),
    .B(_02214_),
    .Y(_02228_)
  );
  OAI21X1 _08868_ (
    .A(_03188_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02229_)
  );
  OAI22X1 _08869_ (
    .A(_03002_),
    .B(_02213_),
    .C(_02228_),
    .D(_02229_),
    .Y(_02050_)
  );
  NOR2X1 _08870_ (
    .A(execution_unit_0.register_file_0.r15_7_ ),
    .B(_02214_),
    .Y(_02230_)
  );
  OAI21X1 _08871_ (
    .A(_03208_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02231_)
  );
  OAI22X1 _08872_ (
    .A(_03004_),
    .B(_02213_),
    .C(_02230_),
    .D(_02231_),
    .Y(_02051_)
  );
  OAI21X1 _08873_ (
    .A(_03227_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02232_)
  );
  INVX1 _08874_ (
    .A(_02232_),
    .Y(_02233_)
  );
  OAI21X1 _08875_ (
    .A(execution_unit_0.register_file_0.r15_8_ ),
    .B(_02214_),
    .C(_02233_),
    .Y(_02234_)
  );
  OAI21X1 _08876_ (
    .A(_03211_),
    .B(_02213_),
    .C(_02234_),
    .Y(_02052_)
  );
  OAI21X1 _08877_ (
    .A(_03244_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02235_)
  );
  INVX1 _08878_ (
    .A(_02235_),
    .Y(_02236_)
  );
  OAI21X1 _08879_ (
    .A(execution_unit_0.register_file_0.r15_9_ ),
    .B(_02214_),
    .C(_02236_),
    .Y(_02237_)
  );
  OAI21X1 _08880_ (
    .A(_03231_),
    .B(_02213_),
    .C(_02237_),
    .Y(_02053_)
  );
  AOI21X1 _08881_ (
    .A(_03265_),
    .B(_02214_),
    .C(_02212_),
    .Y(_02238_)
  );
  OAI21X1 _08882_ (
    .A(execution_unit_0.register_file_0.r15_10_ ),
    .B(_02214_),
    .C(_02238_),
    .Y(_02239_)
  );
  OAI21X1 _08883_ (
    .A(_03248_),
    .B(_02213_),
    .C(_02239_),
    .Y(_02039_)
  );
  OAI21X1 _08884_ (
    .A(_03284_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02240_)
  );
  INVX1 _08885_ (
    .A(_02240_),
    .Y(_02241_)
  );
  OAI21X1 _08886_ (
    .A(execution_unit_0.register_file_0.r15_11_ ),
    .B(_02214_),
    .C(_02241_),
    .Y(_02242_)
  );
  OAI21X1 _08887_ (
    .A(_03268_),
    .B(_02213_),
    .C(_02242_),
    .Y(_02040_)
  );
  OAI21X1 _08888_ (
    .A(execution_unit_0.register_file_0.r15_12_ ),
    .B(_02214_),
    .C(_02213_),
    .Y(_02243_)
  );
  INVX1 _08889_ (
    .A(_02243_),
    .Y(_02244_)
  );
  OAI21X1 _08890_ (
    .A(_03302_),
    .B(_02215_),
    .C(_02244_),
    .Y(_02245_)
  );
  OAI21X1 _08891_ (
    .A(_03288_),
    .B(_02213_),
    .C(_02245_),
    .Y(_02041_)
  );
  OAI21X1 _08892_ (
    .A(execution_unit_0.register_file_0.r15_13_ ),
    .B(_02214_),
    .C(_02213_),
    .Y(_02246_)
  );
  INVX1 _08893_ (
    .A(_02246_),
    .Y(_02247_)
  );
  OAI21X1 _08894_ (
    .A(_03321_),
    .B(_02215_),
    .C(_02247_),
    .Y(_02248_)
  );
  OAI21X1 _08895_ (
    .A(_03306_),
    .B(_02213_),
    .C(_02248_),
    .Y(_02042_)
  );
  OAI21X1 _08896_ (
    .A(execution_unit_0.register_file_0.r15_14_ ),
    .B(_02214_),
    .C(_02213_),
    .Y(_02249_)
  );
  INVX1 _08897_ (
    .A(_02249_),
    .Y(_02250_)
  );
  OAI21X1 _08898_ (
    .A(_02191_),
    .B(_02215_),
    .C(_02250_),
    .Y(_02251_)
  );
  OAI21X1 _08899_ (
    .A(_03325_),
    .B(_02213_),
    .C(_02251_),
    .Y(_02043_)
  );
  OAI21X1 _08900_ (
    .A(execution_unit_0.register_file_0.r15_15_ ),
    .B(_02214_),
    .C(_02213_),
    .Y(_02252_)
  );
  INVX1 _08901_ (
    .A(_02252_),
    .Y(_02253_)
  );
  OAI21X1 _08902_ (
    .A(_02208_),
    .B(_02215_),
    .C(_02253_),
    .Y(_02254_)
  );
  OAI21X1 _08903_ (
    .A(_02195_),
    .B(_02213_),
    .C(_02254_),
    .Y(_02044_)
  );
  AND2X1 _08904_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03031_),
    .Y(_02255_)
  );
  NAND2X1 _08905_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03031_),
    .Y(_02256_)
  );
  AND2X1 _08906_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_1_ ),
    .Y(_02257_)
  );
  NAND2X1 _08907_ (
    .A(execution_unit_0.register_file_0.r1_0_ ),
    .B(_03016_),
    .Y(_02258_)
  );
  OR2X1 _08908_ (
    .A(_02257_),
    .B(_02258_),
    .Y(_02259_)
  );
  NOR2X1 _08909_ (
    .A(_02255_),
    .B(_02259_),
    .Y(_02054_)
  );
  AOI21X1 _08910_ (
    .A(_02985_),
    .B(_02256_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02260_)
  );
  OAI21X1 _08911_ (
    .A(_03093_),
    .B(_02256_),
    .C(_02260_),
    .Y(_02261_)
  );
  AOI21X1 _08912_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_1_ ),
    .C(_02257_),
    .Y(_02262_)
  );
  AOI22X1 _08913_ (
    .A(_02989_),
    .B(_02257_),
    .C(_02261_),
    .D(_02262_),
    .Y(_02061_)
  );
  AOI21X1 _08914_ (
    .A(_03112_),
    .B(_02255_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02263_)
  );
  OAI21X1 _08915_ (
    .A(execution_unit_0.register_file_0.r1_2_ ),
    .B(_02255_),
    .C(_02263_),
    .Y(_02264_)
  );
  AOI21X1 _08916_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_2_ ),
    .C(_02257_),
    .Y(_02265_)
  );
  AOI22X1 _08917_ (
    .A(_02991_),
    .B(_02257_),
    .C(_02264_),
    .D(_02265_),
    .Y(_02062_)
  );
  AOI21X1 _08918_ (
    .A(_02992_),
    .B(_02256_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02266_)
  );
  OAI21X1 _08919_ (
    .A(_03135_),
    .B(_02256_),
    .C(_02266_),
    .Y(_02267_)
  );
  AOI21X1 _08920_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_3_ ),
    .C(_02257_),
    .Y(_02268_)
  );
  AOI22X1 _08921_ (
    .A(_02995_),
    .B(_02257_),
    .C(_02267_),
    .D(_02268_),
    .Y(_02063_)
  );
  AOI21X1 _08922_ (
    .A(_02997_),
    .B(_02256_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02269_)
  );
  OAI21X1 _08923_ (
    .A(_03153_),
    .B(_02256_),
    .C(_02269_),
    .Y(_02270_)
  );
  AOI21X1 _08924_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_4_ ),
    .C(_02257_),
    .Y(_02271_)
  );
  AOI22X1 _08925_ (
    .A(_02998_),
    .B(_02257_),
    .C(_02270_),
    .D(_02271_),
    .Y(_02064_)
  );
  AOI21X1 _08926_ (
    .A(_02999_),
    .B(_02256_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02272_)
  );
  OAI21X1 _08927_ (
    .A(_03171_),
    .B(_02256_),
    .C(_02272_),
    .Y(_02273_)
  );
  AOI21X1 _08928_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_5_ ),
    .C(_02257_),
    .Y(_02274_)
  );
  AOI22X1 _08929_ (
    .A(_03000_),
    .B(_02257_),
    .C(_02273_),
    .D(_02274_),
    .Y(_02065_)
  );
  AOI21X1 _08930_ (
    .A(_03001_),
    .B(_02256_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02275_)
  );
  OAI21X1 _08931_ (
    .A(_03188_),
    .B(_02256_),
    .C(_02275_),
    .Y(_02276_)
  );
  AOI21X1 _08932_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_6_ ),
    .C(_02257_),
    .Y(_02277_)
  );
  AOI22X1 _08933_ (
    .A(_03002_),
    .B(_02257_),
    .C(_02276_),
    .D(_02277_),
    .Y(_02066_)
  );
  AOI21X1 _08934_ (
    .A(_03003_),
    .B(_02256_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02278_)
  );
  OAI21X1 _08935_ (
    .A(_03208_),
    .B(_02256_),
    .C(_02278_),
    .Y(_02279_)
  );
  AOI21X1 _08936_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_7_ ),
    .C(_02257_),
    .Y(_02280_)
  );
  AOI22X1 _08937_ (
    .A(_03004_),
    .B(_02257_),
    .C(_02279_),
    .D(_02280_),
    .Y(_02067_)
  );
  AOI21X1 _08938_ (
    .A(_03005_),
    .B(_02256_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02281_)
  );
  OAI21X1 _08939_ (
    .A(_03227_),
    .B(_02256_),
    .C(_02281_),
    .Y(_02282_)
  );
  AOI21X1 _08940_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_8_ ),
    .C(_02257_),
    .Y(_02283_)
  );
  AOI22X1 _08941_ (
    .A(_03211_),
    .B(_02257_),
    .C(_02282_),
    .D(_02283_),
    .Y(_02068_)
  );
  AOI21X1 _08942_ (
    .A(_03006_),
    .B(_02256_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02284_)
  );
  OAI21X1 _08943_ (
    .A(_03244_),
    .B(_02256_),
    .C(_02284_),
    .Y(_02285_)
  );
  AOI21X1 _08944_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_9_ ),
    .C(_02257_),
    .Y(_02286_)
  );
  AOI22X1 _08945_ (
    .A(_03231_),
    .B(_02257_),
    .C(_02285_),
    .D(_02286_),
    .Y(_02069_)
  );
  AOI21X1 _08946_ (
    .A(_03265_),
    .B(_02255_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02287_)
  );
  OAI21X1 _08947_ (
    .A(execution_unit_0.register_file_0.r1_10_ ),
    .B(_02255_),
    .C(_02287_),
    .Y(_02288_)
  );
  AOI21X1 _08948_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_10_ ),
    .C(_02257_),
    .Y(_02289_)
  );
  AOI22X1 _08949_ (
    .A(_03248_),
    .B(_02257_),
    .C(_02288_),
    .D(_02289_),
    .Y(_02055_)
  );
  AOI21X1 _08950_ (
    .A(_03009_),
    .B(_02256_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02290_)
  );
  OAI21X1 _08951_ (
    .A(_03284_),
    .B(_02256_),
    .C(_02290_),
    .Y(_02291_)
  );
  AOI21X1 _08952_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_11_ ),
    .C(_02257_),
    .Y(_02292_)
  );
  AOI22X1 _08953_ (
    .A(_03268_),
    .B(_02257_),
    .C(_02291_),
    .D(_02292_),
    .Y(_02056_)
  );
  AOI21X1 _08954_ (
    .A(_03010_),
    .B(_02256_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02293_)
  );
  OAI21X1 _08955_ (
    .A(_03302_),
    .B(_02256_),
    .C(_02293_),
    .Y(_02294_)
  );
  AOI21X1 _08956_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_12_ ),
    .C(_02257_),
    .Y(_02295_)
  );
  AOI22X1 _08957_ (
    .A(_03288_),
    .B(_02257_),
    .C(_02294_),
    .D(_02295_),
    .Y(_02057_)
  );
  AOI21X1 _08958_ (
    .A(_03011_),
    .B(_02256_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02296_)
  );
  OAI21X1 _08959_ (
    .A(_03321_),
    .B(_02256_),
    .C(_02296_),
    .Y(_02297_)
  );
  AOI21X1 _08960_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_13_ ),
    .C(_02257_),
    .Y(_02298_)
  );
  AOI22X1 _08961_ (
    .A(_03306_),
    .B(_02257_),
    .C(_02297_),
    .D(_02298_),
    .Y(_02058_)
  );
  AOI21X1 _08962_ (
    .A(_03012_),
    .B(_02256_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02299_)
  );
  OAI21X1 _08963_ (
    .A(_02191_),
    .B(_02256_),
    .C(_02299_),
    .Y(_02300_)
  );
  AOI21X1 _08964_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_14_ ),
    .C(_02257_),
    .Y(_02301_)
  );
  AOI22X1 _08965_ (
    .A(_03325_),
    .B(_02257_),
    .C(_02300_),
    .D(_02301_),
    .Y(_02059_)
  );
  AOI21X1 _08966_ (
    .A(_03015_),
    .B(_02256_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02302_)
  );
  OAI21X1 _08967_ (
    .A(_02208_),
    .B(_02256_),
    .C(_02302_),
    .Y(_02303_)
  );
  AOI21X1 _08968_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_15_ ),
    .C(_02257_),
    .Y(_02304_)
  );
  AOI22X1 _08969_ (
    .A(_02195_),
    .B(_02257_),
    .C(_02303_),
    .D(_02304_),
    .Y(_02060_)
  );
  AOI21X1 _08970_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_2_ ),
    .C(execution_unit_0.reg_sr_wr ),
    .Y(_02305_)
  );
  MUX2X1 _08971_ (
    .A(execution_unit_0.alu_0.status_0_ ),
    .B(execution_unit_0.alu_0.alu_out_0_ ),
    .S(_02305_),
    .Y(_02306_)
  );
  OAI21X1 _08972_ (
    .A(execution_unit_0.alu_0.alu_stat_0_ ),
    .B(_03017_),
    .C(_02980_),
    .Y(_02307_)
  );
  AOI21X1 _08973_ (
    .A(_03017_),
    .B(_02306_),
    .C(_02307_),
    .Y(_02070_)
  );
  MUX2X1 _08974_ (
    .A(execution_unit_0.alu_0.status_1_ ),
    .B(execution_unit_0.alu_0.alu_out_1_ ),
    .S(_02305_),
    .Y(_02308_)
  );
  OAI21X1 _08975_ (
    .A(execution_unit_0.alu_0.Z ),
    .B(_03018_),
    .C(_02980_),
    .Y(_02309_)
  );
  AOI21X1 _08976_ (
    .A(_03018_),
    .B(_02308_),
    .C(_02309_),
    .Y(_02071_)
  );
  MUX2X1 _08977_ (
    .A(execution_unit_0.alu_0.status_2_ ),
    .B(execution_unit_0.alu_0.alu_out_2_ ),
    .S(_02305_),
    .Y(_02310_)
  );
  OAI21X1 _08978_ (
    .A(execution_unit_0.alu_0.N ),
    .B(_03019_),
    .C(_02980_),
    .Y(_02311_)
  );
  AOI21X1 _08979_ (
    .A(_03019_),
    .B(_02310_),
    .C(_02311_),
    .Y(_02072_)
  );
  MUX2X1 _08980_ (
    .A(execution_unit_0.gie ),
    .B(execution_unit_0.alu_0.alu_out_3_ ),
    .S(_02305_),
    .Y(_02312_)
  );
  NOR2X1 _08981_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(_02312_),
    .Y(_02073_)
  );
  OAI21X1 _08982_ (
    .A(_02998_),
    .B(_02305_),
    .C(_02996_),
    .Y(clock_module_0.UNUSED_cpuoff )
  );
  MUX2X1 _08983_ (
    .A(execution_unit_0.register_file_0.r2_4_ ),
    .B(execution_unit_0.alu_0.alu_out_4_ ),
    .S(_02305_),
    .Y(_02313_)
  );
  NOR2X1 _08984_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(_02313_),
    .Y(_02074_)
  );
  MUX2X1 _08985_ (
    .A(clock_module_0.oscoff ),
    .B(execution_unit_0.alu_0.alu_out_5_ ),
    .S(_02305_),
    .Y(_02314_)
  );
  NOR2X1 _08986_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(_02314_),
    .Y(_02075_)
  );
  MUX2X1 _08987_ (
    .A(clock_module_0.scg1 ),
    .B(execution_unit_0.alu_0.alu_out_7_ ),
    .S(_02305_),
    .Y(_02315_)
  );
  NOR2X1 _08988_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(_02315_),
    .Y(_02076_)
  );
  OAI21X1 _08989_ (
    .A(_03211_),
    .B(_02305_),
    .C(_03020_),
    .Y(_02316_)
  );
  AOI21X1 _08990_ (
    .A(execution_unit_0.alu_0.status_3_ ),
    .B(_02305_),
    .C(_02316_),
    .Y(_02317_)
  );
  OAI21X1 _08991_ (
    .A(execution_unit_0.alu_0.alu_stat_3_ ),
    .B(_03020_),
    .C(_02980_),
    .Y(_02318_)
  );
  NOR2X1 _08992_ (
    .A(_02317_),
    .B(_02318_),
    .Y(_02077_)
  );
  AND2X1 _08993_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_4_ ),
    .Y(_02319_)
  );
  NAND2X1 _08994_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_4_ ),
    .Y(_02320_)
  );
  AND2X1 _08995_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03041_),
    .Y(_02321_)
  );
  NAND2X1 _08996_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03041_),
    .Y(_02322_)
  );
  AOI21X1 _08997_ (
    .A(_03069_),
    .B(_02321_),
    .C(_02319_),
    .Y(_02323_)
  );
  OAI21X1 _08998_ (
    .A(execution_unit_0.register_file_0.r4_0_ ),
    .B(_02321_),
    .C(_02323_),
    .Y(_02324_)
  );
  OAI21X1 _08999_ (
    .A(_02984_),
    .B(_02320_),
    .C(_02324_),
    .Y(_02094_)
  );
  AOI21X1 _09000_ (
    .A(_02986_),
    .B(_02322_),
    .C(_02319_),
    .Y(_02325_)
  );
  OAI21X1 _09001_ (
    .A(_03093_),
    .B(_02322_),
    .C(_02325_),
    .Y(_02326_)
  );
  OAI21X1 _09002_ (
    .A(_02989_),
    .B(_02320_),
    .C(_02326_),
    .Y(_02101_)
  );
  AOI21X1 _09003_ (
    .A(_03112_),
    .B(_02321_),
    .C(_02319_),
    .Y(_02327_)
  );
  OAI21X1 _09004_ (
    .A(execution_unit_0.register_file_0.r4_2_ ),
    .B(_02321_),
    .C(_02327_),
    .Y(_02328_)
  );
  OAI21X1 _09005_ (
    .A(_02991_),
    .B(_02320_),
    .C(_02328_),
    .Y(_02102_)
  );
  NOR2X1 _09006_ (
    .A(_03135_),
    .B(_02322_),
    .Y(_02329_)
  );
  OAI21X1 _09007_ (
    .A(execution_unit_0.register_file_0.r4_3_ ),
    .B(_02321_),
    .C(_02320_),
    .Y(_02330_)
  );
  OAI22X1 _09008_ (
    .A(_02995_),
    .B(_02320_),
    .C(_02329_),
    .D(_02330_),
    .Y(_02103_)
  );
  NOR2X1 _09009_ (
    .A(execution_unit_0.register_file_0.r4_4_ ),
    .B(_02321_),
    .Y(_02331_)
  );
  OAI21X1 _09010_ (
    .A(_03153_),
    .B(_02322_),
    .C(_02320_),
    .Y(_02332_)
  );
  OAI22X1 _09011_ (
    .A(_02998_),
    .B(_02320_),
    .C(_02331_),
    .D(_02332_),
    .Y(_02104_)
  );
  NOR2X1 _09012_ (
    .A(execution_unit_0.register_file_0.r4_5_ ),
    .B(_02321_),
    .Y(_02333_)
  );
  OAI21X1 _09013_ (
    .A(_03171_),
    .B(_02322_),
    .C(_02320_),
    .Y(_02334_)
  );
  OAI22X1 _09014_ (
    .A(_03000_),
    .B(_02320_),
    .C(_02333_),
    .D(_02334_),
    .Y(_02105_)
  );
  NOR2X1 _09015_ (
    .A(execution_unit_0.register_file_0.r4_6_ ),
    .B(_02321_),
    .Y(_02335_)
  );
  OAI21X1 _09016_ (
    .A(_03188_),
    .B(_02322_),
    .C(_02320_),
    .Y(_02336_)
  );
  OAI22X1 _09017_ (
    .A(_03002_),
    .B(_02320_),
    .C(_02335_),
    .D(_02336_),
    .Y(_02106_)
  );
  NOR2X1 _09018_ (
    .A(execution_unit_0.register_file_0.r4_7_ ),
    .B(_02321_),
    .Y(_02337_)
  );
  OAI21X1 _09019_ (
    .A(_03208_),
    .B(_02322_),
    .C(_02320_),
    .Y(_02338_)
  );
  OAI22X1 _09020_ (
    .A(_03004_),
    .B(_02320_),
    .C(_02337_),
    .D(_02338_),
    .Y(_02107_)
  );
  OAI21X1 _09021_ (
    .A(_03227_),
    .B(_02322_),
    .C(_02320_),
    .Y(_02339_)
  );
  INVX1 _09022_ (
    .A(_02339_),
    .Y(_02340_)
  );
  OAI21X1 _09023_ (
    .A(execution_unit_0.register_file_0.r4_8_ ),
    .B(_02321_),
    .C(_02340_),
    .Y(_02341_)
  );
  OAI21X1 _09024_ (
    .A(_03211_),
    .B(_02320_),
    .C(_02341_),
    .Y(_02108_)
  );
  OAI21X1 _09025_ (
    .A(_03244_),
    .B(_02322_),
    .C(_02320_),
    .Y(_02342_)
  );
  INVX1 _09026_ (
    .A(_02342_),
    .Y(_02343_)
  );
  OAI21X1 _09027_ (
    .A(execution_unit_0.register_file_0.r4_9_ ),
    .B(_02321_),
    .C(_02343_),
    .Y(_02344_)
  );
  OAI21X1 _09028_ (
    .A(_03231_),
    .B(_02320_),
    .C(_02344_),
    .Y(_02109_)
  );
  AOI21X1 _09029_ (
    .A(_03265_),
    .B(_02321_),
    .C(_02319_),
    .Y(_02345_)
  );
  OAI21X1 _09030_ (
    .A(execution_unit_0.register_file_0.r4_10_ ),
    .B(_02321_),
    .C(_02345_),
    .Y(_02346_)
  );
  OAI21X1 _09031_ (
    .A(_03248_),
    .B(_02320_),
    .C(_02346_),
    .Y(_02095_)
  );
  OAI21X1 _09032_ (
    .A(_03284_),
    .B(_02322_),
    .C(_02320_),
    .Y(_02347_)
  );
  INVX1 _09033_ (
    .A(_02347_),
    .Y(_02348_)
  );
  OAI21X1 _09034_ (
    .A(execution_unit_0.register_file_0.r4_11_ ),
    .B(_02321_),
    .C(_02348_),
    .Y(_02349_)
  );
  OAI21X1 _09035_ (
    .A(_03268_),
    .B(_02320_),
    .C(_02349_),
    .Y(_02096_)
  );
  OAI21X1 _09036_ (
    .A(execution_unit_0.register_file_0.r4_12_ ),
    .B(_02321_),
    .C(_02320_),
    .Y(_02350_)
  );
  INVX1 _09037_ (
    .A(_02350_),
    .Y(_02351_)
  );
  OAI21X1 _09038_ (
    .A(_03302_),
    .B(_02322_),
    .C(_02351_),
    .Y(_02352_)
  );
  OAI21X1 _09039_ (
    .A(_03288_),
    .B(_02320_),
    .C(_02352_),
    .Y(_02097_)
  );
  OAI21X1 _09040_ (
    .A(execution_unit_0.register_file_0.r4_13_ ),
    .B(_02321_),
    .C(_02320_),
    .Y(_02353_)
  );
  INVX1 _09041_ (
    .A(_02353_),
    .Y(_02354_)
  );
  OAI21X1 _09042_ (
    .A(_03321_),
    .B(_02322_),
    .C(_02354_),
    .Y(_02355_)
  );
  OAI21X1 _09043_ (
    .A(_03306_),
    .B(_02320_),
    .C(_02355_),
    .Y(_02098_)
  );
  OAI21X1 _09044_ (
    .A(execution_unit_0.register_file_0.r4_14_ ),
    .B(_02321_),
    .C(_02320_),
    .Y(_02356_)
  );
  INVX1 _09045_ (
    .A(_02356_),
    .Y(_02357_)
  );
  OAI21X1 _09046_ (
    .A(_02191_),
    .B(_02322_),
    .C(_02357_),
    .Y(_02358_)
  );
  OAI21X1 _09047_ (
    .A(_03325_),
    .B(_02320_),
    .C(_02358_),
    .Y(_02099_)
  );
  OAI21X1 _09048_ (
    .A(execution_unit_0.register_file_0.r4_15_ ),
    .B(_02321_),
    .C(_02320_),
    .Y(_02359_)
  );
  INVX1 _09049_ (
    .A(_02359_),
    .Y(_02360_)
  );
  OAI21X1 _09050_ (
    .A(_02208_),
    .B(_02322_),
    .C(_02360_),
    .Y(_02361_)
  );
  OAI21X1 _09051_ (
    .A(_02195_),
    .B(_02320_),
    .C(_02361_),
    .Y(_02100_)
  );
  AND2X1 _09052_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_5_ ),
    .Y(_02362_)
  );
  NAND2X1 _09053_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_5_ ),
    .Y(_02363_)
  );
  AND2X1 _09054_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03054_),
    .Y(_02364_)
  );
  NAND2X1 _09055_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03054_),
    .Y(_02365_)
  );
  AOI21X1 _09056_ (
    .A(_03069_),
    .B(_02364_),
    .C(_02362_),
    .Y(_02366_)
  );
  OAI21X1 _09057_ (
    .A(execution_unit_0.register_file_0.r5_0_ ),
    .B(_02364_),
    .C(_02366_),
    .Y(_02367_)
  );
  OAI21X1 _09058_ (
    .A(_02984_),
    .B(_02363_),
    .C(_02367_),
    .Y(_02110_)
  );
  NOR2X1 _09059_ (
    .A(execution_unit_0.register_file_0.r5_1_ ),
    .B(_02364_),
    .Y(_02368_)
  );
  OAI21X1 _09060_ (
    .A(_03093_),
    .B(_02365_),
    .C(_02363_),
    .Y(_02369_)
  );
  OAI22X1 _09061_ (
    .A(_02989_),
    .B(_02363_),
    .C(_02368_),
    .D(_02369_),
    .Y(_02117_)
  );
  AOI21X1 _09062_ (
    .A(_03112_),
    .B(_02364_),
    .C(_02362_),
    .Y(_02370_)
  );
  OAI21X1 _09063_ (
    .A(execution_unit_0.register_file_0.r5_2_ ),
    .B(_02364_),
    .C(_02370_),
    .Y(_02371_)
  );
  OAI21X1 _09064_ (
    .A(_02991_),
    .B(_02363_),
    .C(_02371_),
    .Y(_02118_)
  );
  NOR2X1 _09065_ (
    .A(execution_unit_0.register_file_0.r5_3_ ),
    .B(_02364_),
    .Y(_02372_)
  );
  OAI21X1 _09066_ (
    .A(_03135_),
    .B(_02365_),
    .C(_02363_),
    .Y(_02373_)
  );
  OAI22X1 _09067_ (
    .A(_02995_),
    .B(_02363_),
    .C(_02372_),
    .D(_02373_),
    .Y(_02119_)
  );
  NOR2X1 _09068_ (
    .A(execution_unit_0.register_file_0.r5_4_ ),
    .B(_02364_),
    .Y(_02374_)
  );
  OAI21X1 _09069_ (
    .A(_03153_),
    .B(_02365_),
    .C(_02363_),
    .Y(_02375_)
  );
  OAI22X1 _09070_ (
    .A(_02998_),
    .B(_02363_),
    .C(_02374_),
    .D(_02375_),
    .Y(_02120_)
  );
  NOR2X1 _09071_ (
    .A(execution_unit_0.register_file_0.r5_5_ ),
    .B(_02364_),
    .Y(_02376_)
  );
  OAI21X1 _09072_ (
    .A(_03171_),
    .B(_02365_),
    .C(_02363_),
    .Y(_02377_)
  );
  OAI22X1 _09073_ (
    .A(_03000_),
    .B(_02363_),
    .C(_02376_),
    .D(_02377_),
    .Y(_02121_)
  );
  NOR2X1 _09074_ (
    .A(execution_unit_0.register_file_0.r5_6_ ),
    .B(_02364_),
    .Y(_02378_)
  );
  OAI21X1 _09075_ (
    .A(_03188_),
    .B(_02365_),
    .C(_02363_),
    .Y(_02379_)
  );
  OAI22X1 _09076_ (
    .A(_03002_),
    .B(_02363_),
    .C(_02378_),
    .D(_02379_),
    .Y(_02122_)
  );
  NOR2X1 _09077_ (
    .A(execution_unit_0.register_file_0.r5_7_ ),
    .B(_02364_),
    .Y(_02380_)
  );
  OAI21X1 _09078_ (
    .A(_03208_),
    .B(_02365_),
    .C(_02363_),
    .Y(_02381_)
  );
  OAI22X1 _09079_ (
    .A(_03004_),
    .B(_02363_),
    .C(_02380_),
    .D(_02381_),
    .Y(_02123_)
  );
  OAI21X1 _09080_ (
    .A(_03227_),
    .B(_02365_),
    .C(_02363_),
    .Y(_02382_)
  );
  INVX1 _09081_ (
    .A(_02382_),
    .Y(_02383_)
  );
  OAI21X1 _09082_ (
    .A(execution_unit_0.register_file_0.r5_8_ ),
    .B(_02364_),
    .C(_02383_),
    .Y(_02384_)
  );
  OAI21X1 _09083_ (
    .A(_03211_),
    .B(_02363_),
    .C(_02384_),
    .Y(_02124_)
  );
  OAI21X1 _09084_ (
    .A(_03244_),
    .B(_02365_),
    .C(_02363_),
    .Y(_02385_)
  );
  INVX1 _09085_ (
    .A(_02385_),
    .Y(_02386_)
  );
  OAI21X1 _09086_ (
    .A(execution_unit_0.register_file_0.r5_9_ ),
    .B(_02364_),
    .C(_02386_),
    .Y(_02387_)
  );
  OAI21X1 _09087_ (
    .A(_03231_),
    .B(_02363_),
    .C(_02387_),
    .Y(_02125_)
  );
  AOI21X1 _09088_ (
    .A(_03265_),
    .B(_02364_),
    .C(_02362_),
    .Y(_02388_)
  );
  OAI21X1 _09089_ (
    .A(execution_unit_0.register_file_0.r5_10_ ),
    .B(_02364_),
    .C(_02388_),
    .Y(_02389_)
  );
  OAI21X1 _09090_ (
    .A(_03248_),
    .B(_02363_),
    .C(_02389_),
    .Y(_02111_)
  );
  OAI21X1 _09091_ (
    .A(_03284_),
    .B(_02365_),
    .C(_02363_),
    .Y(_02390_)
  );
  INVX1 _09092_ (
    .A(_02390_),
    .Y(_02391_)
  );
  OAI21X1 _09093_ (
    .A(execution_unit_0.register_file_0.r5_11_ ),
    .B(_02364_),
    .C(_02391_),
    .Y(_02392_)
  );
  OAI21X1 _09094_ (
    .A(_03268_),
    .B(_02363_),
    .C(_02392_),
    .Y(_02112_)
  );
  OAI21X1 _09095_ (
    .A(execution_unit_0.register_file_0.r5_12_ ),
    .B(_02364_),
    .C(_02363_),
    .Y(_02393_)
  );
  INVX1 _09096_ (
    .A(_02393_),
    .Y(_02394_)
  );
  OAI21X1 _09097_ (
    .A(_03302_),
    .B(_02365_),
    .C(_02394_),
    .Y(_02395_)
  );
  OAI21X1 _09098_ (
    .A(_03288_),
    .B(_02363_),
    .C(_02395_),
    .Y(_02113_)
  );
  OAI21X1 _09099_ (
    .A(execution_unit_0.register_file_0.r5_13_ ),
    .B(_02364_),
    .C(_02363_),
    .Y(_02396_)
  );
  INVX1 _09100_ (
    .A(_02396_),
    .Y(_02397_)
  );
  OAI21X1 _09101_ (
    .A(_03321_),
    .B(_02365_),
    .C(_02397_),
    .Y(_02398_)
  );
  OAI21X1 _09102_ (
    .A(_03306_),
    .B(_02363_),
    .C(_02398_),
    .Y(_02114_)
  );
  OAI21X1 _09103_ (
    .A(execution_unit_0.register_file_0.r5_14_ ),
    .B(_02364_),
    .C(_02363_),
    .Y(_02399_)
  );
  INVX1 _09104_ (
    .A(_02399_),
    .Y(_02400_)
  );
  OAI21X1 _09105_ (
    .A(_02191_),
    .B(_02365_),
    .C(_02400_),
    .Y(_02401_)
  );
  OAI21X1 _09106_ (
    .A(_03325_),
    .B(_02363_),
    .C(_02401_),
    .Y(_02115_)
  );
  OAI21X1 _09107_ (
    .A(execution_unit_0.register_file_0.r5_15_ ),
    .B(_02364_),
    .C(_02363_),
    .Y(_02402_)
  );
  INVX1 _09108_ (
    .A(_02402_),
    .Y(_02403_)
  );
  OAI21X1 _09109_ (
    .A(_02208_),
    .B(_02365_),
    .C(_02403_),
    .Y(_02404_)
  );
  OAI21X1 _09110_ (
    .A(_02195_),
    .B(_02363_),
    .C(_02404_),
    .Y(_02116_)
  );
  NAND2X1 _09111_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_3_ ),
    .Y(_02405_)
  );
  NAND2X1 _09112_ (
    .A(execution_unit_0.register_file_0.r3_0_ ),
    .B(_02405_),
    .Y(_02406_)
  );
  OAI21X1 _09113_ (
    .A(_02984_),
    .B(_02405_),
    .C(_02406_),
    .Y(_02078_)
  );
  NAND2X1 _09114_ (
    .A(execution_unit_0.register_file_0.r3_1_ ),
    .B(_02405_),
    .Y(_02407_)
  );
  OAI21X1 _09115_ (
    .A(_02989_),
    .B(_02405_),
    .C(_02407_),
    .Y(_02085_)
  );
  NAND2X1 _09116_ (
    .A(execution_unit_0.register_file_0.r3_2_ ),
    .B(_02405_),
    .Y(_02408_)
  );
  OAI21X1 _09117_ (
    .A(_02991_),
    .B(_02405_),
    .C(_02408_),
    .Y(_02086_)
  );
  NAND2X1 _09118_ (
    .A(execution_unit_0.register_file_0.r3_3_ ),
    .B(_02405_),
    .Y(_02409_)
  );
  OAI21X1 _09119_ (
    .A(_02995_),
    .B(_02405_),
    .C(_02409_),
    .Y(_02087_)
  );
  NAND2X1 _09120_ (
    .A(execution_unit_0.register_file_0.r3_4_ ),
    .B(_02405_),
    .Y(_02410_)
  );
  OAI21X1 _09121_ (
    .A(_02998_),
    .B(_02405_),
    .C(_02410_),
    .Y(_02088_)
  );
  NAND2X1 _09122_ (
    .A(execution_unit_0.register_file_0.r3_5_ ),
    .B(_02405_),
    .Y(_02411_)
  );
  OAI21X1 _09123_ (
    .A(_03000_),
    .B(_02405_),
    .C(_02411_),
    .Y(_02089_)
  );
  NAND2X1 _09124_ (
    .A(execution_unit_0.register_file_0.r3_6_ ),
    .B(_02405_),
    .Y(_02412_)
  );
  OAI21X1 _09125_ (
    .A(_03002_),
    .B(_02405_),
    .C(_02412_),
    .Y(_02090_)
  );
  NAND2X1 _09126_ (
    .A(execution_unit_0.register_file_0.r3_7_ ),
    .B(_02405_),
    .Y(_02413_)
  );
  OAI21X1 _09127_ (
    .A(_03004_),
    .B(_02405_),
    .C(_02413_),
    .Y(_02091_)
  );
  NAND2X1 _09128_ (
    .A(execution_unit_0.register_file_0.r3_8_ ),
    .B(_02405_),
    .Y(_02414_)
  );
  OAI21X1 _09129_ (
    .A(_03211_),
    .B(_02405_),
    .C(_02414_),
    .Y(_02092_)
  );
  NAND2X1 _09130_ (
    .A(execution_unit_0.register_file_0.r3_9_ ),
    .B(_02405_),
    .Y(_02415_)
  );
  OAI21X1 _09131_ (
    .A(_03231_),
    .B(_02405_),
    .C(_02415_),
    .Y(_02093_)
  );
  NAND2X1 _09132_ (
    .A(execution_unit_0.register_file_0.r3_10_ ),
    .B(_02405_),
    .Y(_02416_)
  );
  OAI21X1 _09133_ (
    .A(_03248_),
    .B(_02405_),
    .C(_02416_),
    .Y(_02079_)
  );
  NAND2X1 _09134_ (
    .A(execution_unit_0.register_file_0.r3_11_ ),
    .B(_02405_),
    .Y(_02417_)
  );
  OAI21X1 _09135_ (
    .A(_03268_),
    .B(_02405_),
    .C(_02417_),
    .Y(_02080_)
  );
  NAND2X1 _09136_ (
    .A(execution_unit_0.register_file_0.r3_12_ ),
    .B(_02405_),
    .Y(_02418_)
  );
  OAI21X1 _09137_ (
    .A(_03288_),
    .B(_02405_),
    .C(_02418_),
    .Y(_02081_)
  );
  NAND2X1 _09138_ (
    .A(execution_unit_0.register_file_0.r3_13_ ),
    .B(_02405_),
    .Y(_02419_)
  );
  OAI21X1 _09139_ (
    .A(_03306_),
    .B(_02405_),
    .C(_02419_),
    .Y(_02082_)
  );
  NAND2X1 _09140_ (
    .A(execution_unit_0.register_file_0.r3_14_ ),
    .B(_02405_),
    .Y(_02420_)
  );
  OAI21X1 _09141_ (
    .A(_03325_),
    .B(_02405_),
    .C(_02420_),
    .Y(_02083_)
  );
  NAND2X1 _09142_ (
    .A(execution_unit_0.register_file_0.r3_15_ ),
    .B(_02405_),
    .Y(_02421_)
  );
  OAI21X1 _09143_ (
    .A(_02195_),
    .B(_02405_),
    .C(_02421_),
    .Y(_02084_)
  );
  AND2X1 _09144_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_6_ ),
    .Y(_02422_)
  );
  NAND2X1 _09145_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_6_ ),
    .Y(_02423_)
  );
  AND2X1 _09146_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03021_),
    .Y(_02424_)
  );
  NAND2X1 _09147_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03021_),
    .Y(_02425_)
  );
  AOI21X1 _09148_ (
    .A(_03069_),
    .B(_02424_),
    .C(_02422_),
    .Y(_02426_)
  );
  OAI21X1 _09149_ (
    .A(execution_unit_0.register_file_0.r6_0_ ),
    .B(_02424_),
    .C(_02426_),
    .Y(_02427_)
  );
  OAI21X1 _09150_ (
    .A(_02984_),
    .B(_02423_),
    .C(_02427_),
    .Y(_02126_)
  );
  NOR2X1 _09151_ (
    .A(execution_unit_0.register_file_0.r6_1_ ),
    .B(_02424_),
    .Y(_02428_)
  );
  OAI21X1 _09152_ (
    .A(_03093_),
    .B(_02425_),
    .C(_02423_),
    .Y(_02429_)
  );
  OAI22X1 _09153_ (
    .A(_02989_),
    .B(_02423_),
    .C(_02428_),
    .D(_02429_),
    .Y(_02133_)
  );
  AOI21X1 _09154_ (
    .A(_03112_),
    .B(_02424_),
    .C(_02422_),
    .Y(_02430_)
  );
  OAI21X1 _09155_ (
    .A(execution_unit_0.register_file_0.r6_2_ ),
    .B(_02424_),
    .C(_02430_),
    .Y(_02431_)
  );
  OAI21X1 _09156_ (
    .A(_02991_),
    .B(_02423_),
    .C(_02431_),
    .Y(_02134_)
  );
  NOR2X1 _09157_ (
    .A(execution_unit_0.register_file_0.r6_3_ ),
    .B(_02424_),
    .Y(_02432_)
  );
  OAI21X1 _09158_ (
    .A(_03135_),
    .B(_02425_),
    .C(_02423_),
    .Y(_02433_)
  );
  OAI22X1 _09159_ (
    .A(_02995_),
    .B(_02423_),
    .C(_02432_),
    .D(_02433_),
    .Y(_02135_)
  );
  NOR2X1 _09160_ (
    .A(execution_unit_0.register_file_0.r6_4_ ),
    .B(_02424_),
    .Y(_02434_)
  );
  OAI21X1 _09161_ (
    .A(_03153_),
    .B(_02425_),
    .C(_02423_),
    .Y(_02435_)
  );
  OAI22X1 _09162_ (
    .A(_02998_),
    .B(_02423_),
    .C(_02434_),
    .D(_02435_),
    .Y(_02136_)
  );
  NOR2X1 _09163_ (
    .A(execution_unit_0.register_file_0.r6_5_ ),
    .B(_02424_),
    .Y(_02436_)
  );
  OAI21X1 _09164_ (
    .A(_03171_),
    .B(_02425_),
    .C(_02423_),
    .Y(_02437_)
  );
  OAI22X1 _09165_ (
    .A(_03000_),
    .B(_02423_),
    .C(_02436_),
    .D(_02437_),
    .Y(_02137_)
  );
  NOR2X1 _09166_ (
    .A(execution_unit_0.register_file_0.r6_6_ ),
    .B(_02424_),
    .Y(_02438_)
  );
  OAI21X1 _09167_ (
    .A(_03188_),
    .B(_02425_),
    .C(_02423_),
    .Y(_02439_)
  );
  OAI22X1 _09168_ (
    .A(_03002_),
    .B(_02423_),
    .C(_02438_),
    .D(_02439_),
    .Y(_02138_)
  );
  NOR2X1 _09169_ (
    .A(execution_unit_0.register_file_0.r6_7_ ),
    .B(_02424_),
    .Y(_02440_)
  );
  OAI21X1 _09170_ (
    .A(_03208_),
    .B(_02425_),
    .C(_02423_),
    .Y(_02441_)
  );
  OAI22X1 _09171_ (
    .A(_03004_),
    .B(_02423_),
    .C(_02440_),
    .D(_02441_),
    .Y(_02139_)
  );
  OAI21X1 _09172_ (
    .A(_03227_),
    .B(_02425_),
    .C(_02423_),
    .Y(_02442_)
  );
  INVX1 _09173_ (
    .A(_02442_),
    .Y(_02443_)
  );
  OAI21X1 _09174_ (
    .A(execution_unit_0.register_file_0.r6_8_ ),
    .B(_02424_),
    .C(_02443_),
    .Y(_02444_)
  );
  OAI21X1 _09175_ (
    .A(_03211_),
    .B(_02423_),
    .C(_02444_),
    .Y(_02140_)
  );
  OAI21X1 _09176_ (
    .A(_03244_),
    .B(_02425_),
    .C(_02423_),
    .Y(_02445_)
  );
  INVX1 _09177_ (
    .A(_02445_),
    .Y(_02446_)
  );
  OAI21X1 _09178_ (
    .A(execution_unit_0.register_file_0.r6_9_ ),
    .B(_02424_),
    .C(_02446_),
    .Y(_02447_)
  );
  OAI21X1 _09179_ (
    .A(_03231_),
    .B(_02423_),
    .C(_02447_),
    .Y(_02141_)
  );
  AOI21X1 _09180_ (
    .A(_03265_),
    .B(_02424_),
    .C(_02422_),
    .Y(_02448_)
  );
  OAI21X1 _09181_ (
    .A(execution_unit_0.register_file_0.r6_10_ ),
    .B(_02424_),
    .C(_02448_),
    .Y(_02449_)
  );
  OAI21X1 _09182_ (
    .A(_03248_),
    .B(_02423_),
    .C(_02449_),
    .Y(_02127_)
  );
  OAI21X1 _09183_ (
    .A(_03284_),
    .B(_02425_),
    .C(_02423_),
    .Y(_02450_)
  );
  INVX1 _09184_ (
    .A(_02450_),
    .Y(_02451_)
  );
  OAI21X1 _09185_ (
    .A(execution_unit_0.register_file_0.r6_11_ ),
    .B(_02424_),
    .C(_02451_),
    .Y(_02452_)
  );
  OAI21X1 _09186_ (
    .A(_03268_),
    .B(_02423_),
    .C(_02452_),
    .Y(_02128_)
  );
  OAI21X1 _09187_ (
    .A(execution_unit_0.register_file_0.r6_12_ ),
    .B(_02424_),
    .C(_02423_),
    .Y(_02453_)
  );
  INVX1 _09188_ (
    .A(_02453_),
    .Y(_02454_)
  );
  OAI21X1 _09189_ (
    .A(_03302_),
    .B(_02425_),
    .C(_02454_),
    .Y(_02455_)
  );
  OAI21X1 _09190_ (
    .A(_03288_),
    .B(_02423_),
    .C(_02455_),
    .Y(_02129_)
  );
  OAI21X1 _09191_ (
    .A(execution_unit_0.register_file_0.r6_13_ ),
    .B(_02424_),
    .C(_02423_),
    .Y(_02456_)
  );
  INVX1 _09192_ (
    .A(_02456_),
    .Y(_02457_)
  );
  OAI21X1 _09193_ (
    .A(_03321_),
    .B(_02425_),
    .C(_02457_),
    .Y(_02458_)
  );
  OAI21X1 _09194_ (
    .A(_03306_),
    .B(_02423_),
    .C(_02458_),
    .Y(_02130_)
  );
  OAI21X1 _09195_ (
    .A(execution_unit_0.register_file_0.r6_14_ ),
    .B(_02424_),
    .C(_02423_),
    .Y(_02459_)
  );
  INVX1 _09196_ (
    .A(_02459_),
    .Y(_02460_)
  );
  OAI21X1 _09197_ (
    .A(_02191_),
    .B(_02425_),
    .C(_02460_),
    .Y(_02461_)
  );
  OAI21X1 _09198_ (
    .A(_03325_),
    .B(_02423_),
    .C(_02461_),
    .Y(_02131_)
  );
  OAI21X1 _09199_ (
    .A(execution_unit_0.register_file_0.r6_15_ ),
    .B(_02424_),
    .C(_02423_),
    .Y(_02462_)
  );
  INVX1 _09200_ (
    .A(_02462_),
    .Y(_02463_)
  );
  OAI21X1 _09201_ (
    .A(_02208_),
    .B(_02425_),
    .C(_02463_),
    .Y(_02464_)
  );
  OAI21X1 _09202_ (
    .A(_02195_),
    .B(_02423_),
    .C(_02464_),
    .Y(_02132_)
  );
  AND2X1 _09203_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_7_ ),
    .Y(_02465_)
  );
  NAND2X1 _09204_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_7_ ),
    .Y(_02466_)
  );
  AND2X1 _09205_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03047_),
    .Y(_02467_)
  );
  NAND2X1 _09206_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03047_),
    .Y(_02468_)
  );
  AOI21X1 _09207_ (
    .A(_03069_),
    .B(_02467_),
    .C(_02465_),
    .Y(_02469_)
  );
  OAI21X1 _09208_ (
    .A(execution_unit_0.register_file_0.r7_0_ ),
    .B(_02467_),
    .C(_02469_),
    .Y(_02470_)
  );
  OAI21X1 _09209_ (
    .A(_02984_),
    .B(_02466_),
    .C(_02470_),
    .Y(_02142_)
  );
  NOR2X1 _09210_ (
    .A(execution_unit_0.register_file_0.r7_1_ ),
    .B(_02467_),
    .Y(_02471_)
  );
  OAI21X1 _09211_ (
    .A(_03093_),
    .B(_02468_),
    .C(_02466_),
    .Y(_02472_)
  );
  OAI22X1 _09212_ (
    .A(_02989_),
    .B(_02466_),
    .C(_02471_),
    .D(_02472_),
    .Y(_02149_)
  );
  AOI21X1 _09213_ (
    .A(_03112_),
    .B(_02467_),
    .C(_02465_),
    .Y(_02473_)
  );
  OAI21X1 _09214_ (
    .A(execution_unit_0.register_file_0.r7_2_ ),
    .B(_02467_),
    .C(_02473_),
    .Y(_02474_)
  );
  OAI21X1 _09215_ (
    .A(_02991_),
    .B(_02466_),
    .C(_02474_),
    .Y(_02150_)
  );
  NOR2X1 _09216_ (
    .A(execution_unit_0.register_file_0.r7_3_ ),
    .B(_02467_),
    .Y(_02475_)
  );
  OAI21X1 _09217_ (
    .A(_03135_),
    .B(_02468_),
    .C(_02466_),
    .Y(_02476_)
  );
  OAI22X1 _09218_ (
    .A(_02995_),
    .B(_02466_),
    .C(_02475_),
    .D(_02476_),
    .Y(_02151_)
  );
  NOR2X1 _09219_ (
    .A(execution_unit_0.register_file_0.r7_4_ ),
    .B(_02467_),
    .Y(_02477_)
  );
  OAI21X1 _09220_ (
    .A(_03153_),
    .B(_02468_),
    .C(_02466_),
    .Y(_02478_)
  );
  OAI22X1 _09221_ (
    .A(_02998_),
    .B(_02466_),
    .C(_02477_),
    .D(_02478_),
    .Y(_02152_)
  );
  NOR2X1 _09222_ (
    .A(execution_unit_0.register_file_0.r7_5_ ),
    .B(_02467_),
    .Y(_02479_)
  );
  OAI21X1 _09223_ (
    .A(_03171_),
    .B(_02468_),
    .C(_02466_),
    .Y(_02480_)
  );
  OAI22X1 _09224_ (
    .A(_03000_),
    .B(_02466_),
    .C(_02479_),
    .D(_02480_),
    .Y(_02153_)
  );
  NOR2X1 _09225_ (
    .A(execution_unit_0.register_file_0.r7_6_ ),
    .B(_02467_),
    .Y(_02481_)
  );
  OAI21X1 _09226_ (
    .A(_03188_),
    .B(_02468_),
    .C(_02466_),
    .Y(_02482_)
  );
  OAI22X1 _09227_ (
    .A(_03002_),
    .B(_02466_),
    .C(_02481_),
    .D(_02482_),
    .Y(_02154_)
  );
  NOR2X1 _09228_ (
    .A(execution_unit_0.register_file_0.r7_7_ ),
    .B(_02467_),
    .Y(_02483_)
  );
  OAI21X1 _09229_ (
    .A(_03208_),
    .B(_02468_),
    .C(_02466_),
    .Y(_02484_)
  );
  OAI22X1 _09230_ (
    .A(_03004_),
    .B(_02466_),
    .C(_02483_),
    .D(_02484_),
    .Y(_02155_)
  );
  OAI21X1 _09231_ (
    .A(_03227_),
    .B(_02468_),
    .C(_02466_),
    .Y(_02485_)
  );
  INVX1 _09232_ (
    .A(_02485_),
    .Y(_02486_)
  );
  OAI21X1 _09233_ (
    .A(execution_unit_0.register_file_0.r7_8_ ),
    .B(_02467_),
    .C(_02486_),
    .Y(_02487_)
  );
  OAI21X1 _09234_ (
    .A(_03211_),
    .B(_02466_),
    .C(_02487_),
    .Y(_02156_)
  );
  OAI21X1 _09235_ (
    .A(_03244_),
    .B(_02468_),
    .C(_02466_),
    .Y(_02488_)
  );
  INVX1 _09236_ (
    .A(_02488_),
    .Y(_02489_)
  );
  OAI21X1 _09237_ (
    .A(execution_unit_0.register_file_0.r7_9_ ),
    .B(_02467_),
    .C(_02489_),
    .Y(_02490_)
  );
  OAI21X1 _09238_ (
    .A(_03231_),
    .B(_02466_),
    .C(_02490_),
    .Y(_02157_)
  );
  OAI21X1 _09239_ (
    .A(execution_unit_0.register_file_0.r7_10_ ),
    .B(_02467_),
    .C(_02466_),
    .Y(_02491_)
  );
  AOI21X1 _09240_ (
    .A(_03265_),
    .B(_02467_),
    .C(_02491_),
    .Y(_02492_)
  );
  INVX1 _09241_ (
    .A(_02492_),
    .Y(_02493_)
  );
  OAI21X1 _09242_ (
    .A(_03248_),
    .B(_02466_),
    .C(_02493_),
    .Y(_02143_)
  );
  OAI21X1 _09243_ (
    .A(_03284_),
    .B(_02468_),
    .C(_02466_),
    .Y(_02494_)
  );
  INVX1 _09244_ (
    .A(_02494_),
    .Y(_02495_)
  );
  OAI21X1 _09245_ (
    .A(execution_unit_0.register_file_0.r7_11_ ),
    .B(_02467_),
    .C(_02495_),
    .Y(_02496_)
  );
  OAI21X1 _09246_ (
    .A(_03268_),
    .B(_02466_),
    .C(_02496_),
    .Y(_02144_)
  );
  OAI21X1 _09247_ (
    .A(execution_unit_0.register_file_0.r7_12_ ),
    .B(_02467_),
    .C(_02466_),
    .Y(_02497_)
  );
  INVX1 _09248_ (
    .A(_02497_),
    .Y(_02498_)
  );
  OAI21X1 _09249_ (
    .A(_03302_),
    .B(_02468_),
    .C(_02498_),
    .Y(_02499_)
  );
  OAI21X1 _09250_ (
    .A(_03288_),
    .B(_02466_),
    .C(_02499_),
    .Y(_02145_)
  );
  OAI21X1 _09251_ (
    .A(execution_unit_0.register_file_0.r7_13_ ),
    .B(_02467_),
    .C(_02466_),
    .Y(_02500_)
  );
  INVX1 _09252_ (
    .A(_02500_),
    .Y(_02501_)
  );
  OAI21X1 _09253_ (
    .A(_03321_),
    .B(_02468_),
    .C(_02501_),
    .Y(_02502_)
  );
  OAI21X1 _09254_ (
    .A(_03306_),
    .B(_02466_),
    .C(_02502_),
    .Y(_02146_)
  );
  OAI21X1 _09255_ (
    .A(execution_unit_0.register_file_0.r7_14_ ),
    .B(_02467_),
    .C(_02466_),
    .Y(_02503_)
  );
  INVX1 _09256_ (
    .A(_02503_),
    .Y(_02504_)
  );
  OAI21X1 _09257_ (
    .A(_02191_),
    .B(_02468_),
    .C(_02504_),
    .Y(_02505_)
  );
  OAI21X1 _09258_ (
    .A(_03325_),
    .B(_02466_),
    .C(_02505_),
    .Y(_02147_)
  );
  OAI21X1 _09259_ (
    .A(execution_unit_0.register_file_0.r7_15_ ),
    .B(_02467_),
    .C(_02466_),
    .Y(_02506_)
  );
  INVX1 _09260_ (
    .A(_02506_),
    .Y(_02507_)
  );
  OAI21X1 _09261_ (
    .A(_02208_),
    .B(_02468_),
    .C(_02507_),
    .Y(_02508_)
  );
  OAI21X1 _09262_ (
    .A(_02195_),
    .B(_02466_),
    .C(_02508_),
    .Y(_02148_)
  );
  AND2X1 _09263_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_8_ ),
    .Y(_02509_)
  );
  NAND2X1 _09264_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_8_ ),
    .Y(_02510_)
  );
  AND2X1 _09265_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03034_),
    .Y(_02511_)
  );
  NAND2X1 _09266_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03034_),
    .Y(_02512_)
  );
  AOI21X1 _09267_ (
    .A(_03069_),
    .B(_02511_),
    .C(_02509_),
    .Y(_02513_)
  );
  OAI21X1 _09268_ (
    .A(execution_unit_0.register_file_0.r8_0_ ),
    .B(_02511_),
    .C(_02513_),
    .Y(_02514_)
  );
  OAI21X1 _09269_ (
    .A(_02984_),
    .B(_02510_),
    .C(_02514_),
    .Y(_02158_)
  );
  NOR2X1 _09270_ (
    .A(execution_unit_0.register_file_0.r8_1_ ),
    .B(_02511_),
    .Y(_02515_)
  );
  OAI21X1 _09271_ (
    .A(_03093_),
    .B(_02512_),
    .C(_02510_),
    .Y(_02516_)
  );
  OAI22X1 _09272_ (
    .A(_02989_),
    .B(_02510_),
    .C(_02515_),
    .D(_02516_),
    .Y(_02165_)
  );
  AOI21X1 _09273_ (
    .A(_03112_),
    .B(_02511_),
    .C(_02509_),
    .Y(_02517_)
  );
  OAI21X1 _09274_ (
    .A(execution_unit_0.register_file_0.r8_2_ ),
    .B(_02511_),
    .C(_02517_),
    .Y(_02518_)
  );
  OAI21X1 _09275_ (
    .A(_02991_),
    .B(_02510_),
    .C(_02518_),
    .Y(_02166_)
  );
  NOR2X1 _09276_ (
    .A(execution_unit_0.register_file_0.r8_3_ ),
    .B(_02511_),
    .Y(_02519_)
  );
  OAI21X1 _09277_ (
    .A(_03135_),
    .B(_02512_),
    .C(_02510_),
    .Y(_02520_)
  );
  OAI22X1 _09278_ (
    .A(_02995_),
    .B(_02510_),
    .C(_02519_),
    .D(_02520_),
    .Y(_02167_)
  );
  NOR2X1 _09279_ (
    .A(execution_unit_0.register_file_0.r8_4_ ),
    .B(_02511_),
    .Y(_02521_)
  );
  OAI21X1 _09280_ (
    .A(_03153_),
    .B(_02512_),
    .C(_02510_),
    .Y(_02522_)
  );
  OAI22X1 _09281_ (
    .A(_02998_),
    .B(_02510_),
    .C(_02521_),
    .D(_02522_),
    .Y(_02168_)
  );
  NOR2X1 _09282_ (
    .A(execution_unit_0.register_file_0.r8_5_ ),
    .B(_02511_),
    .Y(_02523_)
  );
  OAI21X1 _09283_ (
    .A(_03171_),
    .B(_02512_),
    .C(_02510_),
    .Y(_02524_)
  );
  OAI22X1 _09284_ (
    .A(_03000_),
    .B(_02510_),
    .C(_02523_),
    .D(_02524_),
    .Y(_02169_)
  );
  NOR2X1 _09285_ (
    .A(execution_unit_0.register_file_0.r8_6_ ),
    .B(_02511_),
    .Y(_02525_)
  );
  OAI21X1 _09286_ (
    .A(_03188_),
    .B(_02512_),
    .C(_02510_),
    .Y(_02526_)
  );
  OAI22X1 _09287_ (
    .A(_03002_),
    .B(_02510_),
    .C(_02525_),
    .D(_02526_),
    .Y(_02170_)
  );
  NOR2X1 _09288_ (
    .A(execution_unit_0.register_file_0.r8_7_ ),
    .B(_02511_),
    .Y(_02527_)
  );
  OAI21X1 _09289_ (
    .A(_03208_),
    .B(_02512_),
    .C(_02510_),
    .Y(_02528_)
  );
  OAI22X1 _09290_ (
    .A(_03004_),
    .B(_02510_),
    .C(_02527_),
    .D(_02528_),
    .Y(_02171_)
  );
  OAI21X1 _09291_ (
    .A(_03227_),
    .B(_02512_),
    .C(_02510_),
    .Y(_02529_)
  );
  INVX1 _09292_ (
    .A(_02529_),
    .Y(_02530_)
  );
  OAI21X1 _09293_ (
    .A(execution_unit_0.register_file_0.r8_8_ ),
    .B(_02511_),
    .C(_02530_),
    .Y(_02531_)
  );
  OAI21X1 _09294_ (
    .A(_03211_),
    .B(_02510_),
    .C(_02531_),
    .Y(_02172_)
  );
  OAI21X1 _09295_ (
    .A(_03244_),
    .B(_02512_),
    .C(_02510_),
    .Y(_02532_)
  );
  INVX1 _09296_ (
    .A(_02532_),
    .Y(_02533_)
  );
  OAI21X1 _09297_ (
    .A(execution_unit_0.register_file_0.r8_9_ ),
    .B(_02511_),
    .C(_02533_),
    .Y(_02534_)
  );
  OAI21X1 _09298_ (
    .A(_03231_),
    .B(_02510_),
    .C(_02534_),
    .Y(_02173_)
  );
  AOI21X1 _09299_ (
    .A(_03265_),
    .B(_02511_),
    .C(_02509_),
    .Y(_02535_)
  );
  OAI21X1 _09300_ (
    .A(execution_unit_0.register_file_0.r8_10_ ),
    .B(_02511_),
    .C(_02535_),
    .Y(_02536_)
  );
  OAI21X1 _09301_ (
    .A(_03248_),
    .B(_02510_),
    .C(_02536_),
    .Y(_02159_)
  );
  OAI21X1 _09302_ (
    .A(execution_unit_0.register_file_0.r8_11_ ),
    .B(_02511_),
    .C(_02510_),
    .Y(_02537_)
  );
  INVX1 _09303_ (
    .A(_02537_),
    .Y(_02538_)
  );
  OAI21X1 _09304_ (
    .A(_03284_),
    .B(_02512_),
    .C(_02538_),
    .Y(_02539_)
  );
  OAI21X1 _09305_ (
    .A(_03268_),
    .B(_02510_),
    .C(_02539_),
    .Y(_02160_)
  );
  OAI21X1 _09306_ (
    .A(execution_unit_0.register_file_0.r8_12_ ),
    .B(_02511_),
    .C(_02510_),
    .Y(_02540_)
  );
  INVX1 _09307_ (
    .A(_02540_),
    .Y(_02541_)
  );
  OAI21X1 _09308_ (
    .A(_03302_),
    .B(_02512_),
    .C(_02541_),
    .Y(_02542_)
  );
  OAI21X1 _09309_ (
    .A(_03288_),
    .B(_02510_),
    .C(_02542_),
    .Y(_02161_)
  );
  OAI21X1 _09310_ (
    .A(execution_unit_0.register_file_0.r8_13_ ),
    .B(_02511_),
    .C(_02510_),
    .Y(_02543_)
  );
  INVX1 _09311_ (
    .A(_02543_),
    .Y(_02544_)
  );
  OAI21X1 _09312_ (
    .A(_03321_),
    .B(_02512_),
    .C(_02544_),
    .Y(_02545_)
  );
  OAI21X1 _09313_ (
    .A(_03306_),
    .B(_02510_),
    .C(_02545_),
    .Y(_02162_)
  );
  OAI21X1 _09314_ (
    .A(execution_unit_0.register_file_0.r8_14_ ),
    .B(_02511_),
    .C(_02510_),
    .Y(_02546_)
  );
  INVX1 _09315_ (
    .A(_02546_),
    .Y(_02547_)
  );
  OAI21X1 _09316_ (
    .A(_02191_),
    .B(_02512_),
    .C(_02547_),
    .Y(_02548_)
  );
  OAI21X1 _09317_ (
    .A(_03325_),
    .B(_02510_),
    .C(_02548_),
    .Y(_02163_)
  );
  OAI21X1 _09318_ (
    .A(execution_unit_0.register_file_0.r8_15_ ),
    .B(_02511_),
    .C(_02510_),
    .Y(_02549_)
  );
  INVX1 _09319_ (
    .A(_02549_),
    .Y(_02550_)
  );
  OAI21X1 _09320_ (
    .A(_02208_),
    .B(_02512_),
    .C(_02550_),
    .Y(_02551_)
  );
  OAI21X1 _09321_ (
    .A(_02195_),
    .B(_02510_),
    .C(_02551_),
    .Y(_02164_)
  );
  AND2X1 _09322_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_9_ ),
    .Y(_02552_)
  );
  NAND2X1 _09323_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_9_ ),
    .Y(_02553_)
  );
  AND2X1 _09324_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03025_),
    .Y(_02554_)
  );
  NAND2X1 _09325_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03025_),
    .Y(_02555_)
  );
  AOI21X1 _09326_ (
    .A(_03069_),
    .B(_02554_),
    .C(_02552_),
    .Y(_02556_)
  );
  OAI21X1 _09327_ (
    .A(execution_unit_0.register_file_0.r9_0_ ),
    .B(_02554_),
    .C(_02556_),
    .Y(_02557_)
  );
  OAI21X1 _09328_ (
    .A(_02984_),
    .B(_02553_),
    .C(_02557_),
    .Y(_02174_)
  );
  NOR2X1 _09329_ (
    .A(execution_unit_0.register_file_0.r9_1_ ),
    .B(_02554_),
    .Y(_02558_)
  );
  OAI21X1 _09330_ (
    .A(_03093_),
    .B(_02555_),
    .C(_02553_),
    .Y(_02559_)
  );
  OAI22X1 _09331_ (
    .A(_02989_),
    .B(_02553_),
    .C(_02558_),
    .D(_02559_),
    .Y(_02181_)
  );
  AND2X1 _09332_ (
    .A(_03112_),
    .B(_02554_),
    .Y(_02560_)
  );
  OAI21X1 _09333_ (
    .A(execution_unit_0.register_file_0.r9_2_ ),
    .B(_02554_),
    .C(_02553_),
    .Y(_02561_)
  );
  OAI22X1 _09334_ (
    .A(_02991_),
    .B(_02553_),
    .C(_02560_),
    .D(_02561_),
    .Y(_02182_)
  );
  NOR2X1 _09335_ (
    .A(execution_unit_0.register_file_0.r9_3_ ),
    .B(_02554_),
    .Y(_02562_)
  );
  OAI21X1 _09336_ (
    .A(_03135_),
    .B(_02555_),
    .C(_02553_),
    .Y(_02563_)
  );
  OAI22X1 _09337_ (
    .A(_02995_),
    .B(_02553_),
    .C(_02562_),
    .D(_02563_),
    .Y(_02183_)
  );
  NOR2X1 _09338_ (
    .A(execution_unit_0.register_file_0.r9_4_ ),
    .B(_02554_),
    .Y(_02564_)
  );
  OAI21X1 _09339_ (
    .A(_03153_),
    .B(_02555_),
    .C(_02553_),
    .Y(_02565_)
  );
  OAI22X1 _09340_ (
    .A(_02998_),
    .B(_02553_),
    .C(_02564_),
    .D(_02565_),
    .Y(_02184_)
  );
  NOR2X1 _09341_ (
    .A(execution_unit_0.register_file_0.r9_5_ ),
    .B(_02554_),
    .Y(_02566_)
  );
  OAI21X1 _09342_ (
    .A(_03171_),
    .B(_02555_),
    .C(_02553_),
    .Y(_02567_)
  );
  OAI22X1 _09343_ (
    .A(_03000_),
    .B(_02553_),
    .C(_02566_),
    .D(_02567_),
    .Y(_02185_)
  );
  NOR2X1 _09344_ (
    .A(execution_unit_0.register_file_0.r9_6_ ),
    .B(_02554_),
    .Y(_02568_)
  );
  OAI21X1 _09345_ (
    .A(_03188_),
    .B(_02555_),
    .C(_02553_),
    .Y(_02569_)
  );
  OAI22X1 _09346_ (
    .A(_03002_),
    .B(_02553_),
    .C(_02568_),
    .D(_02569_),
    .Y(_02186_)
  );
  NOR2X1 _09347_ (
    .A(execution_unit_0.register_file_0.r9_7_ ),
    .B(_02554_),
    .Y(_02570_)
  );
  OAI21X1 _09348_ (
    .A(_03208_),
    .B(_02555_),
    .C(_02553_),
    .Y(_02571_)
  );
  OAI22X1 _09349_ (
    .A(_03004_),
    .B(_02553_),
    .C(_02570_),
    .D(_02571_),
    .Y(_02187_)
  );
  OAI21X1 _09350_ (
    .A(_03227_),
    .B(_02555_),
    .C(_02553_),
    .Y(_02572_)
  );
  INVX1 _09351_ (
    .A(_02572_),
    .Y(_02573_)
  );
  OAI21X1 _09352_ (
    .A(execution_unit_0.register_file_0.r9_8_ ),
    .B(_02554_),
    .C(_02573_),
    .Y(_02574_)
  );
  OAI21X1 _09353_ (
    .A(_03211_),
    .B(_02553_),
    .C(_02574_),
    .Y(_02188_)
  );
  OAI21X1 _09354_ (
    .A(_03244_),
    .B(_02555_),
    .C(_02553_),
    .Y(_02575_)
  );
  INVX1 _09355_ (
    .A(_02575_),
    .Y(_02576_)
  );
  OAI21X1 _09356_ (
    .A(execution_unit_0.register_file_0.r9_9_ ),
    .B(_02554_),
    .C(_02576_),
    .Y(_02577_)
  );
  OAI21X1 _09357_ (
    .A(_03231_),
    .B(_02553_),
    .C(_02577_),
    .Y(_02189_)
  );
  AOI21X1 _09358_ (
    .A(_03265_),
    .B(_02554_),
    .C(_02552_),
    .Y(_02578_)
  );
  OAI21X1 _09359_ (
    .A(execution_unit_0.register_file_0.r9_10_ ),
    .B(_02554_),
    .C(_02578_),
    .Y(_02579_)
  );
  OAI21X1 _09360_ (
    .A(_03248_),
    .B(_02553_),
    .C(_02579_),
    .Y(_02175_)
  );
  OAI21X1 _09361_ (
    .A(_03284_),
    .B(_02555_),
    .C(_02553_),
    .Y(_02580_)
  );
  INVX1 _09362_ (
    .A(_02580_),
    .Y(_02581_)
  );
  OAI21X1 _09363_ (
    .A(execution_unit_0.register_file_0.r9_11_ ),
    .B(_02554_),
    .C(_02581_),
    .Y(_02582_)
  );
  OAI21X1 _09364_ (
    .A(_03268_),
    .B(_02553_),
    .C(_02582_),
    .Y(_02176_)
  );
  OAI21X1 _09365_ (
    .A(execution_unit_0.register_file_0.r9_12_ ),
    .B(_02554_),
    .C(_02553_),
    .Y(_02583_)
  );
  INVX1 _09366_ (
    .A(_02583_),
    .Y(_02584_)
  );
  OAI21X1 _09367_ (
    .A(_03302_),
    .B(_02555_),
    .C(_02584_),
    .Y(_02585_)
  );
  OAI21X1 _09368_ (
    .A(_03288_),
    .B(_02553_),
    .C(_02585_),
    .Y(_02177_)
  );
  OAI21X1 _09369_ (
    .A(execution_unit_0.register_file_0.r9_13_ ),
    .B(_02554_),
    .C(_02553_),
    .Y(_02586_)
  );
  INVX1 _09370_ (
    .A(_02586_),
    .Y(_02587_)
  );
  OAI21X1 _09371_ (
    .A(_03321_),
    .B(_02555_),
    .C(_02587_),
    .Y(_02588_)
  );
  OAI21X1 _09372_ (
    .A(_03306_),
    .B(_02553_),
    .C(_02588_),
    .Y(_02178_)
  );
  OAI21X1 _09373_ (
    .A(execution_unit_0.register_file_0.r9_14_ ),
    .B(_02554_),
    .C(_02553_),
    .Y(_02589_)
  );
  INVX1 _09374_ (
    .A(_02589_),
    .Y(_02590_)
  );
  OAI21X1 _09375_ (
    .A(_02191_),
    .B(_02555_),
    .C(_02590_),
    .Y(_02591_)
  );
  OAI21X1 _09376_ (
    .A(_03325_),
    .B(_02553_),
    .C(_02591_),
    .Y(_02179_)
  );
  OAI21X1 _09377_ (
    .A(execution_unit_0.register_file_0.r9_15_ ),
    .B(_02554_),
    .C(_02553_),
    .Y(_02592_)
  );
  INVX1 _09378_ (
    .A(_02592_),
    .Y(_02593_)
  );
  OAI21X1 _09379_ (
    .A(_02208_),
    .B(_02555_),
    .C(_02593_),
    .Y(_02594_)
  );
  OAI21X1 _09380_ (
    .A(_02195_),
    .B(_02553_),
    .C(_02594_),
    .Y(_02180_)
  );
  AND2X1 _09381_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_10_ ),
    .Y(_02595_)
  );
  NAND2X1 _09382_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_10_ ),
    .Y(_02596_)
  );
  AND2X1 _09383_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03044_),
    .Y(_02597_)
  );
  NAND2X1 _09384_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03044_),
    .Y(_02598_)
  );
  AOI21X1 _09385_ (
    .A(_03069_),
    .B(_02597_),
    .C(_02595_),
    .Y(_02599_)
  );
  OAI21X1 _09386_ (
    .A(execution_unit_0.register_file_0.r10_0_ ),
    .B(_02597_),
    .C(_02599_),
    .Y(_02600_)
  );
  OAI21X1 _09387_ (
    .A(_02984_),
    .B(_02596_),
    .C(_02600_),
    .Y(_01958_)
  );
  AOI21X1 _09388_ (
    .A(_02988_),
    .B(_02598_),
    .C(_02595_),
    .Y(_02601_)
  );
  OAI21X1 _09389_ (
    .A(_03093_),
    .B(_02598_),
    .C(_02601_),
    .Y(_02602_)
  );
  OAI21X1 _09390_ (
    .A(_02989_),
    .B(_02596_),
    .C(_02602_),
    .Y(_01965_)
  );
  AOI21X1 _09391_ (
    .A(_03112_),
    .B(_02597_),
    .C(_02595_),
    .Y(_02603_)
  );
  OAI21X1 _09392_ (
    .A(execution_unit_0.register_file_0.r10_2_ ),
    .B(_02597_),
    .C(_02603_),
    .Y(_02604_)
  );
  OAI21X1 _09393_ (
    .A(_02991_),
    .B(_02596_),
    .C(_02604_),
    .Y(_01966_)
  );
  NOR2X1 _09394_ (
    .A(execution_unit_0.register_file_0.r10_3_ ),
    .B(_02597_),
    .Y(_02605_)
  );
  OAI21X1 _09395_ (
    .A(_03135_),
    .B(_02598_),
    .C(_02596_),
    .Y(_02606_)
  );
  OAI22X1 _09396_ (
    .A(_02995_),
    .B(_02596_),
    .C(_02605_),
    .D(_02606_),
    .Y(_01967_)
  );
  NOR2X1 _09397_ (
    .A(_03153_),
    .B(_02598_),
    .Y(_02607_)
  );
  OAI21X1 _09398_ (
    .A(execution_unit_0.register_file_0.r10_4_ ),
    .B(_02597_),
    .C(_02596_),
    .Y(_02608_)
  );
  OAI22X1 _09399_ (
    .A(_02998_),
    .B(_02596_),
    .C(_02607_),
    .D(_02608_),
    .Y(_01968_)
  );
  NOR2X1 _09400_ (
    .A(execution_unit_0.register_file_0.r10_5_ ),
    .B(_02597_),
    .Y(_02609_)
  );
  OAI21X1 _09401_ (
    .A(_03171_),
    .B(_02598_),
    .C(_02596_),
    .Y(_02610_)
  );
  OAI22X1 _09402_ (
    .A(_03000_),
    .B(_02596_),
    .C(_02609_),
    .D(_02610_),
    .Y(_01969_)
  );
  NOR2X1 _09403_ (
    .A(execution_unit_0.register_file_0.r10_6_ ),
    .B(_02597_),
    .Y(_02611_)
  );
  OAI21X1 _09404_ (
    .A(_03188_),
    .B(_02598_),
    .C(_02596_),
    .Y(_02612_)
  );
  OAI22X1 _09405_ (
    .A(_03002_),
    .B(_02596_),
    .C(_02611_),
    .D(_02612_),
    .Y(_01970_)
  );
  NOR2X1 _09406_ (
    .A(_03208_),
    .B(_02598_),
    .Y(_02613_)
  );
  OAI21X1 _09407_ (
    .A(execution_unit_0.register_file_0.r10_7_ ),
    .B(_02597_),
    .C(_02596_),
    .Y(_02614_)
  );
  OAI22X1 _09408_ (
    .A(_03004_),
    .B(_02596_),
    .C(_02613_),
    .D(_02614_),
    .Y(_01971_)
  );
  OAI21X1 _09409_ (
    .A(_03227_),
    .B(_02598_),
    .C(_02596_),
    .Y(_02615_)
  );
  INVX1 _09410_ (
    .A(_02615_),
    .Y(_02616_)
  );
  OAI21X1 _09411_ (
    .A(execution_unit_0.register_file_0.r10_8_ ),
    .B(_02597_),
    .C(_02616_),
    .Y(_02617_)
  );
  OAI21X1 _09412_ (
    .A(_03211_),
    .B(_02596_),
    .C(_02617_),
    .Y(_01972_)
  );
  OAI21X1 _09413_ (
    .A(_03244_),
    .B(_02598_),
    .C(_02596_),
    .Y(_02618_)
  );
  INVX1 _09414_ (
    .A(_02618_),
    .Y(_02619_)
  );
  OAI21X1 _09415_ (
    .A(execution_unit_0.register_file_0.r10_9_ ),
    .B(_02597_),
    .C(_02619_),
    .Y(_02620_)
  );
  OAI21X1 _09416_ (
    .A(_03231_),
    .B(_02596_),
    .C(_02620_),
    .Y(_01973_)
  );
  AOI21X1 _09417_ (
    .A(_03265_),
    .B(_02597_),
    .C(_02595_),
    .Y(_02621_)
  );
  OAI21X1 _09418_ (
    .A(execution_unit_0.register_file_0.r10_10_ ),
    .B(_02597_),
    .C(_02621_),
    .Y(_02622_)
  );
  OAI21X1 _09419_ (
    .A(_03248_),
    .B(_02596_),
    .C(_02622_),
    .Y(_01959_)
  );
  OAI21X1 _09420_ (
    .A(_03284_),
    .B(_02598_),
    .C(_02596_),
    .Y(_02623_)
  );
  INVX1 _09421_ (
    .A(_02623_),
    .Y(_02624_)
  );
  OAI21X1 _09422_ (
    .A(execution_unit_0.register_file_0.r10_11_ ),
    .B(_02597_),
    .C(_02624_),
    .Y(_02625_)
  );
  OAI21X1 _09423_ (
    .A(_03268_),
    .B(_02596_),
    .C(_02625_),
    .Y(_01960_)
  );
  OAI21X1 _09424_ (
    .A(execution_unit_0.register_file_0.r10_12_ ),
    .B(_02597_),
    .C(_02596_),
    .Y(_02626_)
  );
  INVX1 _09425_ (
    .A(_02626_),
    .Y(_02627_)
  );
  OAI21X1 _09426_ (
    .A(_03302_),
    .B(_02598_),
    .C(_02627_),
    .Y(_02628_)
  );
  OAI21X1 _09427_ (
    .A(_03288_),
    .B(_02596_),
    .C(_02628_),
    .Y(_01961_)
  );
  OAI21X1 _09428_ (
    .A(execution_unit_0.register_file_0.r10_13_ ),
    .B(_02597_),
    .C(_02596_),
    .Y(_02629_)
  );
  INVX1 _09429_ (
    .A(_02629_),
    .Y(_02630_)
  );
  OAI21X1 _09430_ (
    .A(_03321_),
    .B(_02598_),
    .C(_02630_),
    .Y(_02631_)
  );
  OAI21X1 _09431_ (
    .A(_03306_),
    .B(_02596_),
    .C(_02631_),
    .Y(_01962_)
  );
  OAI21X1 _09432_ (
    .A(execution_unit_0.register_file_0.r10_14_ ),
    .B(_02597_),
    .C(_02596_),
    .Y(_02632_)
  );
  INVX1 _09433_ (
    .A(_02632_),
    .Y(_02633_)
  );
  OAI21X1 _09434_ (
    .A(_02191_),
    .B(_02598_),
    .C(_02633_),
    .Y(_02634_)
  );
  OAI21X1 _09435_ (
    .A(_03325_),
    .B(_02596_),
    .C(_02634_),
    .Y(_01963_)
  );
  OAI21X1 _09436_ (
    .A(execution_unit_0.register_file_0.r10_15_ ),
    .B(_02597_),
    .C(_02596_),
    .Y(_02635_)
  );
  INVX1 _09437_ (
    .A(_02635_),
    .Y(_02636_)
  );
  OAI21X1 _09438_ (
    .A(_02208_),
    .B(_02598_),
    .C(_02636_),
    .Y(_02637_)
  );
  OAI21X1 _09439_ (
    .A(_02195_),
    .B(_02596_),
    .C(_02637_),
    .Y(_01964_)
  );
  AND2X1 _09440_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_11_ ),
    .Y(_02638_)
  );
  NAND2X1 _09441_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_11_ ),
    .Y(_02639_)
  );
  AND2X1 _09442_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03023_),
    .Y(_02640_)
  );
  NAND2X1 _09443_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03023_),
    .Y(_02641_)
  );
  AOI21X1 _09444_ (
    .A(_03069_),
    .B(_02640_),
    .C(_02638_),
    .Y(_02642_)
  );
  OAI21X1 _09445_ (
    .A(execution_unit_0.register_file_0.r11_0_ ),
    .B(_02640_),
    .C(_02642_),
    .Y(_02643_)
  );
  OAI21X1 _09446_ (
    .A(_02984_),
    .B(_02639_),
    .C(_02643_),
    .Y(_01974_)
  );
  NOR2X1 _09447_ (
    .A(execution_unit_0.register_file_0.r11_1_ ),
    .B(_02640_),
    .Y(_02644_)
  );
  OAI21X1 _09448_ (
    .A(_03093_),
    .B(_02641_),
    .C(_02639_),
    .Y(_02645_)
  );
  OAI22X1 _09449_ (
    .A(_02989_),
    .B(_02639_),
    .C(_02644_),
    .D(_02645_),
    .Y(_01981_)
  );
  AOI21X1 _09450_ (
    .A(_03112_),
    .B(_02640_),
    .C(_02638_),
    .Y(_02646_)
  );
  OAI21X1 _09451_ (
    .A(execution_unit_0.register_file_0.r11_2_ ),
    .B(_02640_),
    .C(_02646_),
    .Y(_02647_)
  );
  OAI21X1 _09452_ (
    .A(_02991_),
    .B(_02639_),
    .C(_02647_),
    .Y(_01982_)
  );
  NOR2X1 _09453_ (
    .A(execution_unit_0.register_file_0.r11_3_ ),
    .B(_02640_),
    .Y(_02648_)
  );
  OAI21X1 _09454_ (
    .A(_03135_),
    .B(_02641_),
    .C(_02639_),
    .Y(_02649_)
  );
  OAI22X1 _09455_ (
    .A(_02995_),
    .B(_02639_),
    .C(_02648_),
    .D(_02649_),
    .Y(_01983_)
  );
  NOR2X1 _09456_ (
    .A(execution_unit_0.register_file_0.r11_4_ ),
    .B(_02640_),
    .Y(_02650_)
  );
  OAI21X1 _09457_ (
    .A(_03153_),
    .B(_02641_),
    .C(_02639_),
    .Y(_02651_)
  );
  OAI22X1 _09458_ (
    .A(_02998_),
    .B(_02639_),
    .C(_02650_),
    .D(_02651_),
    .Y(_01984_)
  );
  NOR2X1 _09459_ (
    .A(execution_unit_0.register_file_0.r11_5_ ),
    .B(_02640_),
    .Y(_02652_)
  );
  OAI21X1 _09460_ (
    .A(_03171_),
    .B(_02641_),
    .C(_02639_),
    .Y(_02653_)
  );
  OAI22X1 _09461_ (
    .A(_03000_),
    .B(_02639_),
    .C(_02652_),
    .D(_02653_),
    .Y(_01985_)
  );
  NOR2X1 _09462_ (
    .A(execution_unit_0.register_file_0.r11_6_ ),
    .B(_02640_),
    .Y(_02654_)
  );
  OAI21X1 _09463_ (
    .A(_03188_),
    .B(_02641_),
    .C(_02639_),
    .Y(_02655_)
  );
  OAI22X1 _09464_ (
    .A(_03002_),
    .B(_02639_),
    .C(_02654_),
    .D(_02655_),
    .Y(_01986_)
  );
  NOR2X1 _09465_ (
    .A(_03208_),
    .B(_02641_),
    .Y(_02656_)
  );
  OAI21X1 _09466_ (
    .A(execution_unit_0.register_file_0.r11_7_ ),
    .B(_02640_),
    .C(_02639_),
    .Y(_02657_)
  );
  OAI22X1 _09467_ (
    .A(_03004_),
    .B(_02639_),
    .C(_02656_),
    .D(_02657_),
    .Y(_01987_)
  );
  OAI21X1 _09468_ (
    .A(_03227_),
    .B(_02641_),
    .C(_02639_),
    .Y(_02658_)
  );
  INVX1 _09469_ (
    .A(_02658_),
    .Y(_02659_)
  );
  OAI21X1 _09470_ (
    .A(execution_unit_0.register_file_0.r11_8_ ),
    .B(_02640_),
    .C(_02659_),
    .Y(_02660_)
  );
  OAI21X1 _09471_ (
    .A(_03211_),
    .B(_02639_),
    .C(_02660_),
    .Y(_01988_)
  );
  OAI21X1 _09472_ (
    .A(_03244_),
    .B(_02641_),
    .C(_02639_),
    .Y(_02661_)
  );
  INVX1 _09473_ (
    .A(_02661_),
    .Y(_02662_)
  );
  OAI21X1 _09474_ (
    .A(execution_unit_0.register_file_0.r11_9_ ),
    .B(_02640_),
    .C(_02662_),
    .Y(_02663_)
  );
  OAI21X1 _09475_ (
    .A(_03231_),
    .B(_02639_),
    .C(_02663_),
    .Y(_01989_)
  );
  AOI21X1 _09476_ (
    .A(_03265_),
    .B(_02640_),
    .C(_02638_),
    .Y(_02664_)
  );
  OAI21X1 _09477_ (
    .A(execution_unit_0.register_file_0.r11_10_ ),
    .B(_02640_),
    .C(_02664_),
    .Y(_02665_)
  );
  OAI21X1 _09478_ (
    .A(_03248_),
    .B(_02639_),
    .C(_02665_),
    .Y(_01975_)
  );
  OAI21X1 _09479_ (
    .A(_03284_),
    .B(_02641_),
    .C(_02639_),
    .Y(_02666_)
  );
  INVX1 _09480_ (
    .A(_02666_),
    .Y(_02667_)
  );
  OAI21X1 _09481_ (
    .A(execution_unit_0.register_file_0.r11_11_ ),
    .B(_02640_),
    .C(_02667_),
    .Y(_02668_)
  );
  OAI21X1 _09482_ (
    .A(_03268_),
    .B(_02639_),
    .C(_02668_),
    .Y(_01976_)
  );
  OAI21X1 _09483_ (
    .A(execution_unit_0.register_file_0.r11_12_ ),
    .B(_02640_),
    .C(_02639_),
    .Y(_02669_)
  );
  INVX1 _09484_ (
    .A(_02669_),
    .Y(_02670_)
  );
  OAI21X1 _09485_ (
    .A(_03302_),
    .B(_02641_),
    .C(_02670_),
    .Y(_02671_)
  );
  OAI21X1 _09486_ (
    .A(_03288_),
    .B(_02639_),
    .C(_02671_),
    .Y(_01977_)
  );
  OAI21X1 _09487_ (
    .A(execution_unit_0.register_file_0.r11_13_ ),
    .B(_02640_),
    .C(_02639_),
    .Y(_02672_)
  );
  INVX1 _09488_ (
    .A(_02672_),
    .Y(_02673_)
  );
  OAI21X1 _09489_ (
    .A(_03321_),
    .B(_02641_),
    .C(_02673_),
    .Y(_02674_)
  );
  OAI21X1 _09490_ (
    .A(_03306_),
    .B(_02639_),
    .C(_02674_),
    .Y(_01978_)
  );
  OAI21X1 _09491_ (
    .A(execution_unit_0.register_file_0.r11_14_ ),
    .B(_02640_),
    .C(_02639_),
    .Y(_02675_)
  );
  INVX1 _09492_ (
    .A(_02675_),
    .Y(_02676_)
  );
  OAI21X1 _09493_ (
    .A(_02191_),
    .B(_02641_),
    .C(_02676_),
    .Y(_02677_)
  );
  OAI21X1 _09494_ (
    .A(_03325_),
    .B(_02639_),
    .C(_02677_),
    .Y(_01979_)
  );
  OAI21X1 _09495_ (
    .A(execution_unit_0.register_file_0.r11_15_ ),
    .B(_02640_),
    .C(_02639_),
    .Y(_02678_)
  );
  INVX1 _09496_ (
    .A(_02678_),
    .Y(_02679_)
  );
  OAI21X1 _09497_ (
    .A(_02208_),
    .B(_02641_),
    .C(_02679_),
    .Y(_02680_)
  );
  OAI21X1 _09498_ (
    .A(_02195_),
    .B(_02639_),
    .C(_02680_),
    .Y(_01980_)
  );
  AND2X1 _09499_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_12_ ),
    .Y(_02681_)
  );
  NAND2X1 _09500_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_12_ ),
    .Y(_02682_)
  );
  AND2X1 _09501_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03029_),
    .Y(_02683_)
  );
  NAND2X1 _09502_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03029_),
    .Y(_02684_)
  );
  AOI21X1 _09503_ (
    .A(_03069_),
    .B(_02683_),
    .C(_02681_),
    .Y(_02685_)
  );
  OAI21X1 _09504_ (
    .A(execution_unit_0.register_file_0.r12_0_ ),
    .B(_02683_),
    .C(_02685_),
    .Y(_02686_)
  );
  OAI21X1 _09505_ (
    .A(_02984_),
    .B(_02682_),
    .C(_02686_),
    .Y(_01990_)
  );
  NOR2X1 _09506_ (
    .A(execution_unit_0.register_file_0.r12_1_ ),
    .B(_02683_),
    .Y(_02687_)
  );
  OAI21X1 _09507_ (
    .A(_03093_),
    .B(_02684_),
    .C(_02682_),
    .Y(_02688_)
  );
  OAI22X1 _09508_ (
    .A(_02989_),
    .B(_02682_),
    .C(_02687_),
    .D(_02688_),
    .Y(_01997_)
  );
  NAND2X1 _09509_ (
    .A(execution_unit_0.register_file_0.r12_2_ ),
    .B(_02684_),
    .Y(_02689_)
  );
  OAI21X1 _09510_ (
    .A(_03112_),
    .B(_02684_),
    .C(_02689_),
    .Y(_02690_)
  );
  NAND2X1 _09511_ (
    .A(_02682_),
    .B(_02690_),
    .Y(_02691_)
  );
  OAI21X1 _09512_ (
    .A(_02991_),
    .B(_02682_),
    .C(_02691_),
    .Y(_01998_)
  );
  NOR2X1 _09513_ (
    .A(_03135_),
    .B(_02684_),
    .Y(_02692_)
  );
  OAI21X1 _09514_ (
    .A(execution_unit_0.register_file_0.r12_3_ ),
    .B(_02683_),
    .C(_02682_),
    .Y(_02693_)
  );
  OAI22X1 _09515_ (
    .A(_02995_),
    .B(_02682_),
    .C(_02692_),
    .D(_02693_),
    .Y(_01999_)
  );
  NOR2X1 _09516_ (
    .A(execution_unit_0.register_file_0.r12_4_ ),
    .B(_02683_),
    .Y(_02694_)
  );
  OAI21X1 _09517_ (
    .A(_03153_),
    .B(_02684_),
    .C(_02682_),
    .Y(_02695_)
  );
  OAI22X1 _09518_ (
    .A(_02998_),
    .B(_02682_),
    .C(_02694_),
    .D(_02695_),
    .Y(_02000_)
  );
  NOR2X1 _09519_ (
    .A(execution_unit_0.register_file_0.r12_5_ ),
    .B(_02683_),
    .Y(_02696_)
  );
  OAI21X1 _09520_ (
    .A(_03171_),
    .B(_02684_),
    .C(_02682_),
    .Y(_02697_)
  );
  OAI22X1 _09521_ (
    .A(_03000_),
    .B(_02682_),
    .C(_02696_),
    .D(_02697_),
    .Y(_02001_)
  );
  NOR2X1 _09522_ (
    .A(execution_unit_0.register_file_0.r12_6_ ),
    .B(_02683_),
    .Y(_02698_)
  );
  OAI21X1 _09523_ (
    .A(_03188_),
    .B(_02684_),
    .C(_02682_),
    .Y(_02699_)
  );
  OAI22X1 _09524_ (
    .A(_03002_),
    .B(_02682_),
    .C(_02698_),
    .D(_02699_),
    .Y(_02002_)
  );
  NOR2X1 _09525_ (
    .A(execution_unit_0.register_file_0.r12_7_ ),
    .B(_02683_),
    .Y(_02700_)
  );
  OAI21X1 _09526_ (
    .A(_03208_),
    .B(_02684_),
    .C(_02682_),
    .Y(_02701_)
  );
  OAI22X1 _09527_ (
    .A(_03004_),
    .B(_02682_),
    .C(_02700_),
    .D(_02701_),
    .Y(_02003_)
  );
  OAI21X1 _09528_ (
    .A(execution_unit_0.register_file_0.r12_8_ ),
    .B(_02683_),
    .C(_02682_),
    .Y(_02702_)
  );
  INVX1 _09529_ (
    .A(_02702_),
    .Y(_02703_)
  );
  OAI21X1 _09530_ (
    .A(_03227_),
    .B(_02684_),
    .C(_02703_),
    .Y(_02704_)
  );
  OAI21X1 _09531_ (
    .A(_03211_),
    .B(_02682_),
    .C(_02704_),
    .Y(_02004_)
  );
  OAI21X1 _09532_ (
    .A(_03244_),
    .B(_02684_),
    .C(_02682_),
    .Y(_02705_)
  );
  INVX1 _09533_ (
    .A(_02705_),
    .Y(_02706_)
  );
  OAI21X1 _09534_ (
    .A(execution_unit_0.register_file_0.r12_9_ ),
    .B(_02683_),
    .C(_02706_),
    .Y(_02707_)
  );
  OAI21X1 _09535_ (
    .A(_03231_),
    .B(_02682_),
    .C(_02707_),
    .Y(_02005_)
  );
  AOI21X1 _09536_ (
    .A(_03265_),
    .B(_02683_),
    .C(_02681_),
    .Y(_02708_)
  );
  OAI21X1 _09537_ (
    .A(execution_unit_0.register_file_0.r12_10_ ),
    .B(_02683_),
    .C(_02708_),
    .Y(_02709_)
  );
  OAI21X1 _09538_ (
    .A(_03248_),
    .B(_02682_),
    .C(_02709_),
    .Y(_01991_)
  );
  OAI21X1 _09539_ (
    .A(execution_unit_0.register_file_0.r12_11_ ),
    .B(_02683_),
    .C(_02682_),
    .Y(_02710_)
  );
  INVX1 _09540_ (
    .A(_02710_),
    .Y(_02711_)
  );
  OAI21X1 _09541_ (
    .A(_03284_),
    .B(_02684_),
    .C(_02711_),
    .Y(_02712_)
  );
  OAI21X1 _09542_ (
    .A(_03268_),
    .B(_02682_),
    .C(_02712_),
    .Y(_01992_)
  );
  OAI21X1 _09543_ (
    .A(execution_unit_0.register_file_0.r12_12_ ),
    .B(_02683_),
    .C(_02682_),
    .Y(_02713_)
  );
  INVX1 _09544_ (
    .A(_02713_),
    .Y(_02714_)
  );
  OAI21X1 _09545_ (
    .A(_03302_),
    .B(_02684_),
    .C(_02714_),
    .Y(_02715_)
  );
  OAI21X1 _09546_ (
    .A(_03288_),
    .B(_02682_),
    .C(_02715_),
    .Y(_01993_)
  );
  OAI21X1 _09547_ (
    .A(execution_unit_0.register_file_0.r12_13_ ),
    .B(_02683_),
    .C(_02682_),
    .Y(_02716_)
  );
  INVX1 _09548_ (
    .A(_02716_),
    .Y(_02717_)
  );
  OAI21X1 _09549_ (
    .A(_03321_),
    .B(_02684_),
    .C(_02717_),
    .Y(_02718_)
  );
  OAI21X1 _09550_ (
    .A(_03306_),
    .B(_02682_),
    .C(_02718_),
    .Y(_01994_)
  );
  OAI21X1 _09551_ (
    .A(execution_unit_0.register_file_0.r12_14_ ),
    .B(_02683_),
    .C(_02682_),
    .Y(_02719_)
  );
  INVX1 _09552_ (
    .A(_02719_),
    .Y(_02720_)
  );
  OAI21X1 _09553_ (
    .A(_02191_),
    .B(_02684_),
    .C(_02720_),
    .Y(_02721_)
  );
  OAI21X1 _09554_ (
    .A(_03325_),
    .B(_02682_),
    .C(_02721_),
    .Y(_01995_)
  );
  OAI21X1 _09555_ (
    .A(execution_unit_0.register_file_0.r12_15_ ),
    .B(_02683_),
    .C(_02682_),
    .Y(_02722_)
  );
  INVX1 _09556_ (
    .A(_02722_),
    .Y(_02723_)
  );
  OAI21X1 _09557_ (
    .A(_02208_),
    .B(_02684_),
    .C(_02723_),
    .Y(_02724_)
  );
  OAI21X1 _09558_ (
    .A(_02195_),
    .B(_02682_),
    .C(_02724_),
    .Y(_01996_)
  );
  AND2X1 _09559_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_13_ ),
    .Y(_02725_)
  );
  NAND2X1 _09560_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_13_ ),
    .Y(_02726_)
  );
  AND2X1 _09561_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03038_),
    .Y(_02727_)
  );
  NAND2X1 _09562_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03038_),
    .Y(_02728_)
  );
  AOI21X1 _09563_ (
    .A(_03069_),
    .B(_02727_),
    .C(_02725_),
    .Y(_02729_)
  );
  OAI21X1 _09564_ (
    .A(execution_unit_0.register_file_0.r13_0_ ),
    .B(_02727_),
    .C(_02729_),
    .Y(_02730_)
  );
  OAI21X1 _09565_ (
    .A(_02984_),
    .B(_02726_),
    .C(_02730_),
    .Y(_02006_)
  );
  NOR2X1 _09566_ (
    .A(execution_unit_0.register_file_0.r13_1_ ),
    .B(_02727_),
    .Y(_02731_)
  );
  OAI21X1 _09567_ (
    .A(_03093_),
    .B(_02728_),
    .C(_02726_),
    .Y(_02732_)
  );
  OAI22X1 _09568_ (
    .A(_02989_),
    .B(_02726_),
    .C(_02731_),
    .D(_02732_),
    .Y(_02013_)
  );
  AOI21X1 _09569_ (
    .A(_03112_),
    .B(_02727_),
    .C(_02725_),
    .Y(_02733_)
  );
  OAI21X1 _09570_ (
    .A(execution_unit_0.register_file_0.r13_2_ ),
    .B(_02727_),
    .C(_02733_),
    .Y(_02734_)
  );
  OAI21X1 _09571_ (
    .A(_02991_),
    .B(_02726_),
    .C(_02734_),
    .Y(_02014_)
  );
  AOI21X1 _09572_ (
    .A(_02994_),
    .B(_02728_),
    .C(_02725_),
    .Y(_02735_)
  );
  OAI21X1 _09573_ (
    .A(_03135_),
    .B(_02728_),
    .C(_02735_),
    .Y(_02736_)
  );
  OAI21X1 _09574_ (
    .A(_02995_),
    .B(_02726_),
    .C(_02736_),
    .Y(_02015_)
  );
  NOR2X1 _09575_ (
    .A(execution_unit_0.register_file_0.r13_4_ ),
    .B(_02727_),
    .Y(_02737_)
  );
  OAI21X1 _09576_ (
    .A(_03153_),
    .B(_02728_),
    .C(_02726_),
    .Y(_02738_)
  );
  OAI22X1 _09577_ (
    .A(_02998_),
    .B(_02726_),
    .C(_02737_),
    .D(_02738_),
    .Y(_02016_)
  );
  NOR2X1 _09578_ (
    .A(execution_unit_0.register_file_0.r13_5_ ),
    .B(_02727_),
    .Y(_02739_)
  );
  OAI21X1 _09579_ (
    .A(_03171_),
    .B(_02728_),
    .C(_02726_),
    .Y(_02740_)
  );
  OAI22X1 _09580_ (
    .A(_03000_),
    .B(_02726_),
    .C(_02739_),
    .D(_02740_),
    .Y(_02017_)
  );
  NOR2X1 _09581_ (
    .A(execution_unit_0.register_file_0.r13_6_ ),
    .B(_02727_),
    .Y(_02741_)
  );
  OAI21X1 _09582_ (
    .A(_03188_),
    .B(_02728_),
    .C(_02726_),
    .Y(_02742_)
  );
  OAI22X1 _09583_ (
    .A(_03002_),
    .B(_02726_),
    .C(_02741_),
    .D(_02742_),
    .Y(_02018_)
  );
  NOR2X1 _09584_ (
    .A(execution_unit_0.register_file_0.r13_7_ ),
    .B(_02727_),
    .Y(_02743_)
  );
  OAI21X1 _09585_ (
    .A(_03208_),
    .B(_02728_),
    .C(_02726_),
    .Y(_02744_)
  );
  OAI22X1 _09586_ (
    .A(_03004_),
    .B(_02726_),
    .C(_02743_),
    .D(_02744_),
    .Y(_02019_)
  );
  OAI21X1 _09587_ (
    .A(_03227_),
    .B(_02728_),
    .C(_02726_),
    .Y(_02745_)
  );
  INVX1 _09588_ (
    .A(_02745_),
    .Y(_02746_)
  );
  OAI21X1 _09589_ (
    .A(execution_unit_0.register_file_0.r13_8_ ),
    .B(_02727_),
    .C(_02746_),
    .Y(_02747_)
  );
  OAI21X1 _09590_ (
    .A(_03211_),
    .B(_02726_),
    .C(_02747_),
    .Y(_02020_)
  );
  AOI21X1 _09591_ (
    .A(_03007_),
    .B(_02728_),
    .C(_02725_),
    .Y(_02748_)
  );
  OAI21X1 _09592_ (
    .A(_03244_),
    .B(_02728_),
    .C(_02748_),
    .Y(_02749_)
  );
  OAI21X1 _09593_ (
    .A(_03231_),
    .B(_02726_),
    .C(_02749_),
    .Y(_02021_)
  );
  AOI21X1 _09594_ (
    .A(_03265_),
    .B(_02727_),
    .C(_02725_),
    .Y(_02750_)
  );
  OAI21X1 _09595_ (
    .A(execution_unit_0.register_file_0.r13_10_ ),
    .B(_02727_),
    .C(_02750_),
    .Y(_02751_)
  );
  OAI21X1 _09596_ (
    .A(_03248_),
    .B(_02726_),
    .C(_02751_),
    .Y(_02007_)
  );
  OAI21X1 _09597_ (
    .A(_03284_),
    .B(_02728_),
    .C(_02726_),
    .Y(_02752_)
  );
  INVX1 _09598_ (
    .A(_02752_),
    .Y(_02753_)
  );
  OAI21X1 _09599_ (
    .A(execution_unit_0.register_file_0.r13_11_ ),
    .B(_02727_),
    .C(_02753_),
    .Y(_02754_)
  );
  OAI21X1 _09600_ (
    .A(_03268_),
    .B(_02726_),
    .C(_02754_),
    .Y(_02008_)
  );
  OAI21X1 _09601_ (
    .A(execution_unit_0.register_file_0.r13_12_ ),
    .B(_02727_),
    .C(_02726_),
    .Y(_02755_)
  );
  INVX1 _09602_ (
    .A(_02755_),
    .Y(_02756_)
  );
  OAI21X1 _09603_ (
    .A(_03302_),
    .B(_02728_),
    .C(_02756_),
    .Y(_02757_)
  );
  OAI21X1 _09604_ (
    .A(_03288_),
    .B(_02726_),
    .C(_02757_),
    .Y(_02009_)
  );
  OAI21X1 _09605_ (
    .A(execution_unit_0.register_file_0.r13_13_ ),
    .B(_02727_),
    .C(_02726_),
    .Y(_02758_)
  );
  INVX1 _09606_ (
    .A(_02758_),
    .Y(_02759_)
  );
  OAI21X1 _09607_ (
    .A(_03321_),
    .B(_02728_),
    .C(_02759_),
    .Y(_02760_)
  );
  OAI21X1 _09608_ (
    .A(_03306_),
    .B(_02726_),
    .C(_02760_),
    .Y(_02010_)
  );
  OAI21X1 _09609_ (
    .A(execution_unit_0.register_file_0.r13_14_ ),
    .B(_02727_),
    .C(_02726_),
    .Y(_02761_)
  );
  INVX1 _09610_ (
    .A(_02761_),
    .Y(_02762_)
  );
  OAI21X1 _09611_ (
    .A(_02191_),
    .B(_02728_),
    .C(_02762_),
    .Y(_02763_)
  );
  OAI21X1 _09612_ (
    .A(_03325_),
    .B(_02726_),
    .C(_02763_),
    .Y(_02011_)
  );
  OAI21X1 _09613_ (
    .A(execution_unit_0.register_file_0.r13_15_ ),
    .B(_02727_),
    .C(_02726_),
    .Y(_02764_)
  );
  INVX1 _09614_ (
    .A(_02764_),
    .Y(_02765_)
  );
  OAI21X1 _09615_ (
    .A(_02208_),
    .B(_02728_),
    .C(_02765_),
    .Y(_02766_)
  );
  OAI21X1 _09616_ (
    .A(_02195_),
    .B(_02726_),
    .C(_02766_),
    .Y(_02012_)
  );
  AOI21X1 _09617_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_0_ ),
    .C(execution_unit_0.reg_pc_call ),
    .Y(_02767_)
  );
  INVX1 _09618_ (
    .A(_02767_),
    .Y(execution_unit_0.pc_sw_wr )
  );
  AOI22X1 _09619_ (
    .A(execution_unit_0.register_file_0.r14_0_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_0_ ),
    .Y(_02768_)
  );
  AOI22X1 _09620_ (
    .A(execution_unit_0.register_file_0.r10_0_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_0_ ),
    .Y(_02769_)
  );
  NAND2X1 _09621_ (
    .A(_02768_),
    .B(_02769_),
    .Y(_02770_)
  );
  AOI22X1 _09622_ (
    .A(execution_unit_0.register_file_0.r15_0_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .C(execution_unit_0.inst_dest_9_ ),
    .D(execution_unit_0.register_file_0.r9_0_ ),
    .Y(_02771_)
  );
  AOI22X1 _09623_ (
    .A(execution_unit_0.register_file_0.r11_0_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_0_ ),
    .Y(_02772_)
  );
  NAND2X1 _09624_ (
    .A(_02771_),
    .B(_02772_),
    .Y(_02773_)
  );
  NOR2X1 _09625_ (
    .A(_02770_),
    .B(_02773_),
    .Y(_02774_)
  );
  AOI22X1 _09626_ (
    .A(execution_unit_0.register_file_0.r7_0_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_0_ ),
    .Y(_02775_)
  );
  AOI22X1 _09627_ (
    .A(execution_unit_0.register_file_0.r5_0_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_0_ ),
    .Y(_02776_)
  );
  NAND2X1 _09628_ (
    .A(_02775_),
    .B(_02776_),
    .Y(_02777_)
  );
  AOI22X1 _09629_ (
    .A(execution_unit_0.register_file_0.r4_0_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_0_ ),
    .Y(_02778_)
  );
  AOI22X1 _09630_ (
    .A(execution_unit_0.register_file_0.r1_0_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .C(execution_unit_0.inst_dest_2_ ),
    .D(execution_unit_0.alu_0.status_0_ ),
    .Y(_02779_)
  );
  NAND2X1 _09631_ (
    .A(_02778_),
    .B(_02779_),
    .Y(_02780_)
  );
  NOR2X1 _09632_ (
    .A(_02777_),
    .B(_02780_),
    .Y(_02781_)
  );
  NAND2X1 _09633_ (
    .A(_02774_),
    .B(_02781_),
    .Y(dbg_0.dbg_reg_din_0_ )
  );
  AOI22X1 _09634_ (
    .A(execution_unit_0.register_file_0.r15_1_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_1_ ),
    .Y(_02782_)
  );
  AOI22X1 _09635_ (
    .A(execution_unit_0.register_file_0.r4_1_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_1_ ),
    .Y(_02783_)
  );
  NAND2X1 _09636_ (
    .A(_02782_),
    .B(_02783_),
    .Y(_02784_)
  );
  AOI22X1 _09637_ (
    .A(execution_unit_0.register_file_0.r7_1_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .C(execution_unit_0.inst_dest_9_ ),
    .D(execution_unit_0.register_file_0.r9_1_ ),
    .Y(_02785_)
  );
  AOI22X1 _09638_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_1_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_1_ ),
    .Y(_02786_)
  );
  NAND2X1 _09639_ (
    .A(_02785_),
    .B(_02786_),
    .Y(_02787_)
  );
  NOR2X1 _09640_ (
    .A(_02784_),
    .B(_02787_),
    .Y(_02788_)
  );
  AOI22X1 _09641_ (
    .A(execution_unit_0.alu_0.status_1_ ),
    .B(execution_unit_0.inst_dest_2_ ),
    .C(execution_unit_0.inst_dest_10_ ),
    .D(execution_unit_0.register_file_0.r10_1_ ),
    .Y(_02789_)
  );
  AOI22X1 _09642_ (
    .A(execution_unit_0.register_file_0.r13_1_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_1_ ),
    .Y(_02790_)
  );
  NAND2X1 _09643_ (
    .A(_02789_),
    .B(_02790_),
    .Y(_02791_)
  );
  AOI22X1 _09644_ (
    .A(execution_unit_0.register_file_0.r5_1_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_1_ ),
    .Y(_02792_)
  );
  AOI22X1 _09645_ (
    .A(execution_unit_0.register_file_0.r3_1_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_1_ ),
    .Y(_02793_)
  );
  NAND2X1 _09646_ (
    .A(_02792_),
    .B(_02793_),
    .Y(_02794_)
  );
  NOR2X1 _09647_ (
    .A(_02791_),
    .B(_02794_),
    .Y(_02795_)
  );
  NAND2X1 _09648_ (
    .A(_02788_),
    .B(_02795_),
    .Y(dbg_0.dbg_reg_din_1_ )
  );
  AOI22X1 _09649_ (
    .A(execution_unit_0.register_file_0.r15_2_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_2_ ),
    .Y(_02796_)
  );
  AOI22X1 _09650_ (
    .A(execution_unit_0.alu_0.status_2_ ),
    .B(execution_unit_0.inst_dest_2_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_2_ ),
    .Y(_02797_)
  );
  NAND2X1 _09651_ (
    .A(_02796_),
    .B(_02797_),
    .Y(_02798_)
  );
  AOI22X1 _09652_ (
    .A(execution_unit_0.register_file_0.r1_2_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_2_ ),
    .Y(_02799_)
  );
  AOI22X1 _09653_ (
    .A(execution_unit_0.register_file_0.r4_2_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_2_ ),
    .Y(_02800_)
  );
  NAND2X1 _09654_ (
    .A(_02799_),
    .B(_02800_),
    .Y(_02801_)
  );
  NOR2X1 _09655_ (
    .A(_02798_),
    .B(_02801_),
    .Y(_02802_)
  );
  AOI22X1 _09656_ (
    .A(execution_unit_0.register_file_0.r11_2_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_2_ ),
    .Y(_02803_)
  );
  AOI22X1 _09657_ (
    .A(execution_unit_0.register_file_0.r9_2_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_10_ ),
    .D(execution_unit_0.register_file_0.r10_2_ ),
    .Y(_02804_)
  );
  NAND2X1 _09658_ (
    .A(_02803_),
    .B(_02804_),
    .Y(_02805_)
  );
  AOI22X1 _09659_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_2_ ),
    .C(execution_unit_0.register_file_0.r12_2_ ),
    .D(execution_unit_0.inst_dest_12_ ),
    .Y(_02806_)
  );
  AOI22X1 _09660_ (
    .A(execution_unit_0.register_file_0.r5_2_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_2_ ),
    .Y(_02807_)
  );
  NAND2X1 _09661_ (
    .A(_02806_),
    .B(_02807_),
    .Y(_02808_)
  );
  NOR2X1 _09662_ (
    .A(_02805_),
    .B(_02808_),
    .Y(_02809_)
  );
  NAND2X1 _09663_ (
    .A(_02802_),
    .B(_02809_),
    .Y(dbg_0.dbg_reg_din_2_ )
  );
  AOI22X1 _09664_ (
    .A(execution_unit_0.register_file_0.r15_3_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_3_ ),
    .Y(_02810_)
  );
  AOI22X1 _09665_ (
    .A(execution_unit_0.register_file_0.r4_3_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(execution_unit_0.inst_dest_10_ ),
    .D(execution_unit_0.register_file_0.r10_3_ ),
    .Y(_02811_)
  );
  NAND2X1 _09666_ (
    .A(_02810_),
    .B(_02811_),
    .Y(_02812_)
  );
  AOI22X1 _09667_ (
    .A(execution_unit_0.register_file_0.r11_3_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_3_ ),
    .Y(_02813_)
  );
  AOI22X1 _09668_ (
    .A(execution_unit_0.register_file_0.r3_3_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_3_ ),
    .Y(_02814_)
  );
  NAND2X1 _09669_ (
    .A(_02813_),
    .B(_02814_),
    .Y(_02815_)
  );
  NOR2X1 _09670_ (
    .A(_02812_),
    .B(_02815_),
    .Y(_02816_)
  );
  AOI22X1 _09671_ (
    .A(execution_unit_0.register_file_0.r1_3_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_3_ ),
    .Y(_02817_)
  );
  AOI22X1 _09672_ (
    .A(execution_unit_0.gie ),
    .B(execution_unit_0.inst_dest_2_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_3_ ),
    .Y(_02818_)
  );
  NAND2X1 _09673_ (
    .A(_02817_),
    .B(_02818_),
    .Y(_02819_)
  );
  AOI22X1 _09674_ (
    .A(execution_unit_0.register_file_0.r5_3_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_9_ ),
    .D(execution_unit_0.register_file_0.r9_3_ ),
    .Y(_02820_)
  );
  AOI22X1 _09675_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_3_ ),
    .C(execution_unit_0.register_file_0.r13_3_ ),
    .D(execution_unit_0.inst_dest_13_ ),
    .Y(_02821_)
  );
  NAND2X1 _09676_ (
    .A(_02820_),
    .B(_02821_),
    .Y(_02822_)
  );
  NOR2X1 _09677_ (
    .A(_02819_),
    .B(_02822_),
    .Y(_02823_)
  );
  NAND2X1 _09678_ (
    .A(_02816_),
    .B(_02823_),
    .Y(dbg_0.dbg_reg_din_3_ )
  );
  AOI22X1 _09679_ (
    .A(execution_unit_0.register_file_0.r8_4_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_4_ ),
    .Y(_02824_)
  );
  AOI22X1 _09680_ (
    .A(execution_unit_0.register_file_0.r7_4_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_4_ ),
    .Y(_02825_)
  );
  NAND2X1 _09681_ (
    .A(_02824_),
    .B(_02825_),
    .Y(_02826_)
  );
  AOI22X1 _09682_ (
    .A(execution_unit_0.register_file_0.r15_4_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_4_ ),
    .Y(_02827_)
  );
  AOI22X1 _09683_ (
    .A(execution_unit_0.register_file_0.r10_4_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_4_ ),
    .Y(_02828_)
  );
  NAND2X1 _09684_ (
    .A(_02827_),
    .B(_02828_),
    .Y(_02829_)
  );
  NOR2X1 _09685_ (
    .A(_02826_),
    .B(_02829_),
    .Y(_02830_)
  );
  AOI22X1 _09686_ (
    .A(execution_unit_0.register_file_0.r5_4_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_4_ ),
    .Y(_02831_)
  );
  AOI22X1 _09687_ (
    .A(execution_unit_0.register_file_0.r1_4_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .C(execution_unit_0.inst_dest_9_ ),
    .D(execution_unit_0.register_file_0.r9_4_ ),
    .Y(_02832_)
  );
  NAND2X1 _09688_ (
    .A(_02831_),
    .B(_02832_),
    .Y(_02833_)
  );
  AOI22X1 _09689_ (
    .A(execution_unit_0.register_file_0.r2_4_ ),
    .B(execution_unit_0.inst_dest_2_ ),
    .C(execution_unit_0.inst_dest_4_ ),
    .D(execution_unit_0.register_file_0.r4_4_ ),
    .Y(_02834_)
  );
  AOI22X1 _09690_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_4_ ),
    .C(execution_unit_0.register_file_0.r6_4_ ),
    .D(execution_unit_0.inst_dest_6_ ),
    .Y(_02835_)
  );
  NAND2X1 _09691_ (
    .A(_02834_),
    .B(_02835_),
    .Y(_02836_)
  );
  NOR2X1 _09692_ (
    .A(_02833_),
    .B(_02836_),
    .Y(_02837_)
  );
  NAND2X1 _09693_ (
    .A(_02830_),
    .B(_02837_),
    .Y(dbg_0.dbg_reg_din_4_ )
  );
  AOI22X1 _09694_ (
    .A(clock_module_0.oscoff ),
    .B(execution_unit_0.inst_dest_2_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_5_ ),
    .Y(_02838_)
  );
  AOI22X1 _09695_ (
    .A(execution_unit_0.register_file_0.r6_5_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .C(execution_unit_0.inst_dest_9_ ),
    .D(execution_unit_0.register_file_0.r9_5_ ),
    .Y(_02839_)
  );
  NAND2X1 _09696_ (
    .A(_02838_),
    .B(_02839_),
    .Y(_02840_)
  );
  AOI22X1 _09697_ (
    .A(execution_unit_0.register_file_0.r15_5_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_5_ ),
    .Y(_02841_)
  );
  AOI22X1 _09698_ (
    .A(execution_unit_0.register_file_0.r10_5_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_5_ ),
    .Y(_02842_)
  );
  NAND2X1 _09699_ (
    .A(_02841_),
    .B(_02842_),
    .Y(_02843_)
  );
  NOR2X1 _09700_ (
    .A(_02840_),
    .B(_02843_),
    .Y(_02844_)
  );
  AOI22X1 _09701_ (
    .A(execution_unit_0.register_file_0.r5_5_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_5_ ),
    .Y(_02845_)
  );
  AOI22X1 _09702_ (
    .A(execution_unit_0.register_file_0.r7_5_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_5_ ),
    .Y(_02846_)
  );
  NAND2X1 _09703_ (
    .A(_02845_),
    .B(_02846_),
    .Y(_02847_)
  );
  AOI22X1 _09704_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_5_ ),
    .C(execution_unit_0.register_file_0.r4_5_ ),
    .D(execution_unit_0.inst_dest_4_ ),
    .Y(_02848_)
  );
  AOI22X1 _09705_ (
    .A(execution_unit_0.register_file_0.r1_5_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_5_ ),
    .Y(_02849_)
  );
  NAND2X1 _09706_ (
    .A(_02848_),
    .B(_02849_),
    .Y(_02850_)
  );
  NOR2X1 _09707_ (
    .A(_02847_),
    .B(_02850_),
    .Y(_02851_)
  );
  NAND2X1 _09708_ (
    .A(_02844_),
    .B(_02851_),
    .Y(dbg_0.dbg_reg_din_5_ )
  );
  NAND2X1 _09709_ (
    .A(execution_unit_0.register_file_0.r12_6_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .Y(_02852_)
  );
  NAND2X1 _09710_ (
    .A(execution_unit_0.register_file_0.r6_6_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .Y(_02853_)
  );
  AOI22X1 _09711_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_6_ ),
    .C(execution_unit_0.register_file_0.r15_6_ ),
    .D(execution_unit_0.inst_dest_15_ ),
    .Y(_02854_)
  );
  NAND2X1 _09712_ (
    .A(_02852_),
    .B(_02854_),
    .Y(_02855_)
  );
  AOI22X1 _09713_ (
    .A(execution_unit_0.register_file_0.r1_6_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_6_ ),
    .Y(_02856_)
  );
  AOI22X1 _09714_ (
    .A(execution_unit_0.register_file_0.r3_6_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_6_ ),
    .Y(_02857_)
  );
  AOI22X1 _09715_ (
    .A(execution_unit_0.register_file_0.r5_6_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_6_ ),
    .Y(_02858_)
  );
  NAND3X1 _09716_ (
    .A(_02856_),
    .B(_02857_),
    .C(_02858_),
    .Y(_02859_)
  );
  AOI21X1 _09717_ (
    .A(execution_unit_0.register_file_0.r4_6_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(_02859_),
    .Y(_02860_)
  );
  AOI22X1 _09718_ (
    .A(execution_unit_0.register_file_0.r9_6_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_6_ ),
    .Y(_02861_)
  );
  AOI22X1 _09719_ (
    .A(execution_unit_0.register_file_0.r8_6_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(execution_unit_0.inst_dest_10_ ),
    .D(execution_unit_0.register_file_0.r10_6_ ),
    .Y(_02862_)
  );
  NAND2X1 _09720_ (
    .A(_02853_),
    .B(_02862_),
    .Y(_02863_)
  );
  NOR2X1 _09721_ (
    .A(_02855_),
    .B(_02863_),
    .Y(_02864_)
  );
  NAND3X1 _09722_ (
    .A(_02860_),
    .B(_02861_),
    .C(_02864_),
    .Y(dbg_0.dbg_reg_din_6_ )
  );
  AOI22X1 _09723_ (
    .A(execution_unit_0.register_file_0.r15_7_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_7_ ),
    .Y(_02865_)
  );
  AOI22X1 _09724_ (
    .A(execution_unit_0.register_file_0.r6_7_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_7_ ),
    .Y(_02866_)
  );
  NAND2X1 _09725_ (
    .A(_02865_),
    .B(_02866_),
    .Y(_02867_)
  );
  AOI22X1 _09726_ (
    .A(clock_module_0.scg1 ),
    .B(execution_unit_0.inst_dest_2_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_7_ ),
    .Y(_02868_)
  );
  AOI22X1 _09727_ (
    .A(execution_unit_0.register_file_0.r5_7_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_7_ ),
    .Y(_02869_)
  );
  NAND2X1 _09728_ (
    .A(_02868_),
    .B(_02869_),
    .Y(_02870_)
  );
  NOR2X1 _09729_ (
    .A(_02867_),
    .B(_02870_),
    .Y(_02871_)
  );
  AOI22X1 _09730_ (
    .A(execution_unit_0.register_file_0.r12_7_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_7_ ),
    .Y(_02872_)
  );
  AOI22X1 _09731_ (
    .A(execution_unit_0.register_file_0.r9_7_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_10_ ),
    .D(execution_unit_0.register_file_0.r10_7_ ),
    .Y(_02873_)
  );
  NAND2X1 _09732_ (
    .A(_02872_),
    .B(_02873_),
    .Y(_02874_)
  );
  AOI22X1 _09733_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_7_ ),
    .C(execution_unit_0.register_file_0.r4_7_ ),
    .D(execution_unit_0.inst_dest_4_ ),
    .Y(_02875_)
  );
  AOI22X1 _09734_ (
    .A(execution_unit_0.register_file_0.r7_7_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_7_ ),
    .Y(_02876_)
  );
  NAND2X1 _09735_ (
    .A(_02875_),
    .B(_02876_),
    .Y(_02877_)
  );
  NOR2X1 _09736_ (
    .A(_02874_),
    .B(_02877_),
    .Y(_02878_)
  );
  NAND2X1 _09737_ (
    .A(_02871_),
    .B(_02878_),
    .Y(dbg_0.dbg_reg_din_7_ )
  );
  AOI22X1 _09738_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_8_ ),
    .C(execution_unit_0.register_file_0.r5_8_ ),
    .D(execution_unit_0.inst_dest_5_ ),
    .Y(_02879_)
  );
  AOI22X1 _09739_ (
    .A(execution_unit_0.register_file_0.r1_8_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .C(execution_unit_0.inst_dest_9_ ),
    .D(execution_unit_0.register_file_0.r9_8_ ),
    .Y(_02880_)
  );
  NAND2X1 _09740_ (
    .A(_02879_),
    .B(_02880_),
    .Y(_02881_)
  );
  AOI22X1 _09741_ (
    .A(execution_unit_0.register_file_0.r15_8_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_8_ ),
    .Y(_02882_)
  );
  AOI22X1 _09742_ (
    .A(execution_unit_0.alu_0.status_3_ ),
    .B(execution_unit_0.inst_dest_2_ ),
    .C(execution_unit_0.inst_dest_10_ ),
    .D(execution_unit_0.register_file_0.r10_8_ ),
    .Y(_02883_)
  );
  NAND2X1 _09743_ (
    .A(_02882_),
    .B(_02883_),
    .Y(_02884_)
  );
  NOR2X1 _09744_ (
    .A(_02881_),
    .B(_02884_),
    .Y(_02885_)
  );
  AOI22X1 _09745_ (
    .A(execution_unit_0.register_file_0.r3_8_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_8_ ),
    .Y(_02886_)
  );
  AOI22X1 _09746_ (
    .A(execution_unit_0.register_file_0.r12_8_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_8_ ),
    .Y(_02887_)
  );
  NAND2X1 _09747_ (
    .A(_02886_),
    .B(_02887_),
    .Y(_02888_)
  );
  AOI22X1 _09748_ (
    .A(execution_unit_0.register_file_0.r4_8_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_8_ ),
    .Y(_02889_)
  );
  AOI22X1 _09749_ (
    .A(execution_unit_0.register_file_0.r6_8_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_8_ ),
    .Y(_02890_)
  );
  NAND2X1 _09750_ (
    .A(_02889_),
    .B(_02890_),
    .Y(_02891_)
  );
  NOR2X1 _09751_ (
    .A(_02888_),
    .B(_02891_),
    .Y(_02892_)
  );
  NAND2X1 _09752_ (
    .A(_02885_),
    .B(_02892_),
    .Y(dbg_0.dbg_reg_din_8_ )
  );
  NAND2X1 _09753_ (
    .A(execution_unit_0.register_file_0.r10_9_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .Y(_02893_)
  );
  NAND2X1 _09754_ (
    .A(execution_unit_0.register_file_0.r9_9_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .Y(_02894_)
  );
  AOI22X1 _09755_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_9_ ),
    .C(execution_unit_0.register_file_0.r15_9_ ),
    .D(execution_unit_0.inst_dest_15_ ),
    .Y(_02895_)
  );
  NAND2X1 _09756_ (
    .A(_02894_),
    .B(_02895_),
    .Y(_02896_)
  );
  AOI21X1 _09757_ (
    .A(execution_unit_0.register_file_0.r1_9_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .C(_02896_),
    .Y(_02897_)
  );
  AOI22X1 _09758_ (
    .A(execution_unit_0.register_file_0.r11_9_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_9_ ),
    .Y(_02898_)
  );
  AOI22X1 _09759_ (
    .A(execution_unit_0.register_file_0.r3_9_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_9_ ),
    .Y(_02899_)
  );
  NAND2X1 _09760_ (
    .A(_02898_),
    .B(_02899_),
    .Y(_02900_)
  );
  AOI21X1 _09761_ (
    .A(execution_unit_0.register_file_0.r5_9_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(_02900_),
    .Y(_02901_)
  );
  AOI22X1 _09762_ (
    .A(execution_unit_0.register_file_0.r6_9_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_9_ ),
    .Y(_02902_)
  );
  AOI22X1 _09763_ (
    .A(execution_unit_0.register_file_0.r4_9_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_9_ ),
    .Y(_02903_)
  );
  NAND3X1 _09764_ (
    .A(_02893_),
    .B(_02902_),
    .C(_02903_),
    .Y(_02904_)
  );
  AOI21X1 _09765_ (
    .A(execution_unit_0.register_file_0.r8_9_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(_02904_),
    .Y(_02905_)
  );
  NAND3X1 _09766_ (
    .A(_02897_),
    .B(_02901_),
    .C(_02905_),
    .Y(dbg_0.dbg_reg_din_9_ )
  );
  AOI22X1 _09767_ (
    .A(execution_unit_0.register_file_0.r5_10_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_10_ ),
    .Y(_02906_)
  );
  NAND2X1 _09768_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_10_ ),
    .Y(_02907_)
  );
  NAND2X1 _09769_ (
    .A(execution_unit_0.register_file_0.r12_10_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .Y(_02908_)
  );
  AOI22X1 _09770_ (
    .A(execution_unit_0.register_file_0.r15_10_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_10_ ),
    .Y(_02909_)
  );
  NAND2X1 _09771_ (
    .A(_02908_),
    .B(_02909_),
    .Y(_02910_)
  );
  AOI22X1 _09772_ (
    .A(execution_unit_0.register_file_0.r9_10_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_10_ ),
    .Y(_02911_)
  );
  AOI22X1 _09773_ (
    .A(execution_unit_0.register_file_0.r3_10_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_10_ ),
    .Y(_02912_)
  );
  NAND3X1 _09774_ (
    .A(_02906_),
    .B(_02911_),
    .C(_02912_),
    .Y(_02913_)
  );
  AOI21X1 _09775_ (
    .A(execution_unit_0.register_file_0.r4_10_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(_02913_),
    .Y(_02914_)
  );
  AOI22X1 _09776_ (
    .A(execution_unit_0.register_file_0.r1_10_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_10_ ),
    .Y(_02915_)
  );
  AOI22X1 _09777_ (
    .A(execution_unit_0.register_file_0.r8_10_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(execution_unit_0.inst_dest_10_ ),
    .D(execution_unit_0.register_file_0.r10_10_ ),
    .Y(_02916_)
  );
  NAND2X1 _09778_ (
    .A(_02907_),
    .B(_02916_),
    .Y(_02917_)
  );
  NOR2X1 _09779_ (
    .A(_02910_),
    .B(_02917_),
    .Y(_02918_)
  );
  NAND3X1 _09780_ (
    .A(_02914_),
    .B(_02915_),
    .C(_02918_),
    .Y(dbg_0.dbg_reg_din_10_ )
  );
  AOI22X1 _09781_ (
    .A(execution_unit_0.register_file_0.r7_11_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_11_ ),
    .Y(_02919_)
  );
  AOI22X1 _09782_ (
    .A(execution_unit_0.register_file_0.r1_11_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_11_ ),
    .Y(_02920_)
  );
  AND2X1 _09783_ (
    .A(_02919_),
    .B(_02920_),
    .Y(_02921_)
  );
  AOI22X1 _09784_ (
    .A(execution_unit_0.register_file_0.r5_11_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_11_ ),
    .Y(_02922_)
  );
  AOI22X1 _09785_ (
    .A(execution_unit_0.register_file_0.r4_11_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_11_ ),
    .Y(_02923_)
  );
  NAND3X1 _09786_ (
    .A(_02921_),
    .B(_02922_),
    .C(_02923_),
    .Y(_02924_)
  );
  AOI22X1 _09787_ (
    .A(execution_unit_0.register_file_0.r15_11_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_11_ ),
    .Y(_02925_)
  );
  INVX1 _09788_ (
    .A(_02925_),
    .Y(_02926_)
  );
  AOI21X1 _09789_ (
    .A(execution_unit_0.register_file_0.r10_11_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(_02926_),
    .Y(_02927_)
  );
  AOI22X1 _09790_ (
    .A(execution_unit_0.register_file_0.r3_11_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_11_ ),
    .Y(_02928_)
  );
  AOI22X1 _09791_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_11_ ),
    .C(execution_unit_0.inst_dest_9_ ),
    .D(execution_unit_0.register_file_0.r9_11_ ),
    .Y(_02929_)
  );
  NAND3X1 _09792_ (
    .A(_02927_),
    .B(_02928_),
    .C(_02929_),
    .Y(_02930_)
  );
  OR2X1 _09793_ (
    .A(_02924_),
    .B(_02930_),
    .Y(dbg_0.dbg_reg_din_11_ )
  );
  AOI22X1 _09794_ (
    .A(execution_unit_0.register_file_0.r5_12_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_12_ ),
    .Y(_02931_)
  );
  AOI22X1 _09795_ (
    .A(execution_unit_0.register_file_0.r15_12_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_12_ ),
    .Y(_02932_)
  );
  AND2X1 _09796_ (
    .A(_02931_),
    .B(_02932_),
    .Y(_02933_)
  );
  AOI22X1 _09797_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_12_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_12_ ),
    .Y(_02934_)
  );
  AOI22X1 _09798_ (
    .A(execution_unit_0.register_file_0.r4_12_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_12_ ),
    .Y(_02935_)
  );
  NAND3X1 _09799_ (
    .A(_02933_),
    .B(_02934_),
    .C(_02935_),
    .Y(_02936_)
  );
  AOI22X1 _09800_ (
    .A(execution_unit_0.register_file_0.r3_12_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(execution_unit_0.inst_dest_10_ ),
    .D(execution_unit_0.register_file_0.r10_12_ ),
    .Y(_02937_)
  );
  INVX1 _09801_ (
    .A(_02937_),
    .Y(_02938_)
  );
  AOI21X1 _09802_ (
    .A(execution_unit_0.register_file_0.r7_12_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .C(_02938_),
    .Y(_02939_)
  );
  AOI22X1 _09803_ (
    .A(execution_unit_0.register_file_0.r12_12_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_12_ ),
    .Y(_02940_)
  );
  AOI22X1 _09804_ (
    .A(execution_unit_0.register_file_0.r9_12_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_12_ ),
    .Y(_02941_)
  );
  NAND3X1 _09805_ (
    .A(_02939_),
    .B(_02940_),
    .C(_02941_),
    .Y(_02942_)
  );
  OR2X1 _09806_ (
    .A(_02936_),
    .B(_02942_),
    .Y(dbg_0.dbg_reg_din_12_ )
  );
  NAND2X1 _09807_ (
    .A(execution_unit_0.register_file_0.r4_13_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .Y(_02943_)
  );
  NAND2X1 _09808_ (
    .A(execution_unit_0.register_file_0.r15_13_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .Y(_02944_)
  );
  AOI22X1 _09809_ (
    .A(execution_unit_0.register_file_0.r9_13_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_13_ ),
    .Y(_02945_)
  );
  AOI22X1 _09810_ (
    .A(execution_unit_0.register_file_0.r8_13_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(execution_unit_0.inst_dest_10_ ),
    .D(execution_unit_0.register_file_0.r10_13_ ),
    .Y(_02946_)
  );
  AOI22X1 _09811_ (
    .A(execution_unit_0.register_file_0.r6_13_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_13_ ),
    .Y(_02947_)
  );
  NAND2X1 _09812_ (
    .A(_02946_),
    .B(_02947_),
    .Y(_02948_)
  );
  AOI21X1 _09813_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_13_ ),
    .C(_02948_),
    .Y(_02949_)
  );
  NAND3X1 _09814_ (
    .A(_02943_),
    .B(_02944_),
    .C(_02945_),
    .Y(_02950_)
  );
  AOI22X1 _09815_ (
    .A(execution_unit_0.register_file_0.r1_13_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_13_ ),
    .Y(_02951_)
  );
  AOI22X1 _09816_ (
    .A(execution_unit_0.register_file_0.r3_13_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_13_ ),
    .Y(_02952_)
  );
  AOI22X1 _09817_ (
    .A(execution_unit_0.register_file_0.r5_13_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_13_ ),
    .Y(_02953_)
  );
  NAND3X1 _09818_ (
    .A(_02951_),
    .B(_02952_),
    .C(_02953_),
    .Y(_02954_)
  );
  NOR2X1 _09819_ (
    .A(_02950_),
    .B(_02954_),
    .Y(_02955_)
  );
  NAND2X1 _09820_ (
    .A(_02949_),
    .B(_02955_),
    .Y(dbg_0.dbg_reg_din_13_ )
  );
  AOI22X1 _09821_ (
    .A(execution_unit_0.register_file_0.r4_14_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_14_ ),
    .Y(_02956_)
  );
  AOI22X1 _09822_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_14_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_14_ ),
    .Y(_02957_)
  );
  AOI22X1 _09823_ (
    .A(execution_unit_0.register_file_0.r9_14_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_10_ ),
    .D(execution_unit_0.register_file_0.r10_14_ ),
    .Y(_02958_)
  );
  AOI22X1 _09824_ (
    .A(execution_unit_0.register_file_0.r11_14_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_14_ ),
    .Y(_02959_)
  );
  AND2X1 _09825_ (
    .A(_02958_),
    .B(_02959_),
    .Y(_02960_)
  );
  NAND3X1 _09826_ (
    .A(_02956_),
    .B(_02957_),
    .C(_02960_),
    .Y(_02961_)
  );
  AOI22X1 _09827_ (
    .A(execution_unit_0.register_file_0.r5_14_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_14_ ),
    .Y(_02962_)
  );
  INVX1 _09828_ (
    .A(_02962_),
    .Y(_02963_)
  );
  AOI21X1 _09829_ (
    .A(execution_unit_0.register_file_0.r8_14_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(_02963_),
    .Y(_02964_)
  );
  AOI22X1 _09830_ (
    .A(execution_unit_0.register_file_0.r3_14_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_14_ ),
    .Y(_02965_)
  );
  AOI22X1 _09831_ (
    .A(execution_unit_0.register_file_0.r15_14_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_14_ ),
    .Y(_02966_)
  );
  NAND3X1 _09832_ (
    .A(_02964_),
    .B(_02965_),
    .C(_02966_),
    .Y(_02967_)
  );
  OR2X1 _09833_ (
    .A(_02961_),
    .B(_02967_),
    .Y(dbg_0.dbg_reg_din_14_ )
  );
  AOI22X1 _09834_ (
    .A(execution_unit_0.inst_dest_14_ ),
    .B(execution_unit_0.register_file_0.r14_15_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_15_ ),
    .Y(_02968_)
  );
  AOI22X1 _09835_ (
    .A(execution_unit_0.register_file_0.r4_15_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_15_ ),
    .Y(_02969_)
  );
  AND2X1 _09836_ (
    .A(_02968_),
    .B(_02969_),
    .Y(_02970_)
  );
  AOI22X1 _09837_ (
    .A(execution_unit_0.register_file_0.r7_15_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_15_ ),
    .Y(_02971_)
  );
  AOI22X1 _09838_ (
    .A(execution_unit_0.register_file_0.r10_15_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_15_ ),
    .Y(_02972_)
  );
  NAND3X1 _09839_ (
    .A(_02970_),
    .B(_02971_),
    .C(_02972_),
    .Y(_02973_)
  );
  AOI22X1 _09840_ (
    .A(execution_unit_0.register_file_0.r5_15_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_15_ ),
    .Y(_02974_)
  );
  INVX1 _09841_ (
    .A(_02974_),
    .Y(_02975_)
  );
  AOI21X1 _09842_ (
    .A(execution_unit_0.register_file_0.r6_15_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .C(_02975_),
    .Y(_02976_)
  );
  AOI22X1 _09843_ (
    .A(execution_unit_0.register_file_0.r9_15_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_15_ ),
    .Y(_02977_)
  );
  AOI22X1 _09844_ (
    .A(execution_unit_0.register_file_0.r15_15_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_15_ ),
    .Y(_02978_)
  );
  NAND3X1 _09845_ (
    .A(_02976_),
    .B(_02977_),
    .C(_02978_),
    .Y(_02979_)
  );
  OR2X1 _09846_ (
    .A(_02973_),
    .B(_02979_),
    .Y(dbg_0.dbg_reg_din_15_ )
  );
  DFFSR _09847_ (
    .CLK(dco_clk),
    .D(_02038_),
    .Q(execution_unit_0.register_file_0.r15_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09848_ (
    .CLK(dco_clk),
    .D(_02045_),
    .Q(execution_unit_0.register_file_0.r15_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09849_ (
    .CLK(dco_clk),
    .D(_02046_),
    .Q(execution_unit_0.register_file_0.r15_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09850_ (
    .CLK(dco_clk),
    .D(_02047_),
    .Q(execution_unit_0.register_file_0.r15_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09851_ (
    .CLK(dco_clk),
    .D(_02048_),
    .Q(execution_unit_0.register_file_0.r15_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09852_ (
    .CLK(dco_clk),
    .D(_02049_),
    .Q(execution_unit_0.register_file_0.r15_5_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09853_ (
    .CLK(dco_clk),
    .D(_02050_),
    .Q(execution_unit_0.register_file_0.r15_6_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09854_ (
    .CLK(dco_clk),
    .D(_02051_),
    .Q(execution_unit_0.register_file_0.r15_7_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09855_ (
    .CLK(dco_clk),
    .D(_02052_),
    .Q(execution_unit_0.register_file_0.r15_8_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09856_ (
    .CLK(dco_clk),
    .D(_02053_),
    .Q(execution_unit_0.register_file_0.r15_9_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09857_ (
    .CLK(dco_clk),
    .D(_02039_),
    .Q(execution_unit_0.register_file_0.r15_10_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09858_ (
    .CLK(dco_clk),
    .D(_02040_),
    .Q(execution_unit_0.register_file_0.r15_11_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09859_ (
    .CLK(dco_clk),
    .D(_02041_),
    .Q(execution_unit_0.register_file_0.r15_12_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09860_ (
    .CLK(dco_clk),
    .D(_02042_),
    .Q(execution_unit_0.register_file_0.r15_13_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09861_ (
    .CLK(dco_clk),
    .D(_02043_),
    .Q(execution_unit_0.register_file_0.r15_14_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09862_ (
    .CLK(dco_clk),
    .D(_02044_),
    .Q(execution_unit_0.register_file_0.r15_15_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09863_ (
    .CLK(dco_clk),
    .D(_02022_),
    .Q(execution_unit_0.register_file_0.r14_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09864_ (
    .CLK(dco_clk),
    .D(_02029_),
    .Q(execution_unit_0.register_file_0.r14_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09865_ (
    .CLK(dco_clk),
    .D(_02030_),
    .Q(execution_unit_0.register_file_0.r14_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09866_ (
    .CLK(dco_clk),
    .D(_02031_),
    .Q(execution_unit_0.register_file_0.r14_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09867_ (
    .CLK(dco_clk),
    .D(_02032_),
    .Q(execution_unit_0.register_file_0.r14_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09868_ (
    .CLK(dco_clk),
    .D(_02033_),
    .Q(execution_unit_0.register_file_0.r14_5_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09869_ (
    .CLK(dco_clk),
    .D(_02034_),
    .Q(execution_unit_0.register_file_0.r14_6_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09870_ (
    .CLK(dco_clk),
    .D(_02035_),
    .Q(execution_unit_0.register_file_0.r14_7_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09871_ (
    .CLK(dco_clk),
    .D(_02036_),
    .Q(execution_unit_0.register_file_0.r14_8_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09872_ (
    .CLK(dco_clk),
    .D(_02037_),
    .Q(execution_unit_0.register_file_0.r14_9_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09873_ (
    .CLK(dco_clk),
    .D(_02023_),
    .Q(execution_unit_0.register_file_0.r14_10_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09874_ (
    .CLK(dco_clk),
    .D(_02024_),
    .Q(execution_unit_0.register_file_0.r14_11_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09875_ (
    .CLK(dco_clk),
    .D(_02025_),
    .Q(execution_unit_0.register_file_0.r14_12_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09876_ (
    .CLK(dco_clk),
    .D(_02026_),
    .Q(execution_unit_0.register_file_0.r14_13_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09877_ (
    .CLK(dco_clk),
    .D(_02027_),
    .Q(execution_unit_0.register_file_0.r14_14_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09878_ (
    .CLK(dco_clk),
    .D(_02028_),
    .Q(execution_unit_0.register_file_0.r14_15_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09879_ (
    .CLK(dco_clk),
    .D(_02006_),
    .Q(execution_unit_0.register_file_0.r13_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09880_ (
    .CLK(dco_clk),
    .D(_02013_),
    .Q(execution_unit_0.register_file_0.r13_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09881_ (
    .CLK(dco_clk),
    .D(_02014_),
    .Q(execution_unit_0.register_file_0.r13_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09882_ (
    .CLK(dco_clk),
    .D(_02015_),
    .Q(execution_unit_0.register_file_0.r13_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09883_ (
    .CLK(dco_clk),
    .D(_02016_),
    .Q(execution_unit_0.register_file_0.r13_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09884_ (
    .CLK(dco_clk),
    .D(_02017_),
    .Q(execution_unit_0.register_file_0.r13_5_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09885_ (
    .CLK(dco_clk),
    .D(_02018_),
    .Q(execution_unit_0.register_file_0.r13_6_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09886_ (
    .CLK(dco_clk),
    .D(_02019_),
    .Q(execution_unit_0.register_file_0.r13_7_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09887_ (
    .CLK(dco_clk),
    .D(_02020_),
    .Q(execution_unit_0.register_file_0.r13_8_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09888_ (
    .CLK(dco_clk),
    .D(_02021_),
    .Q(execution_unit_0.register_file_0.r13_9_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09889_ (
    .CLK(dco_clk),
    .D(_02007_),
    .Q(execution_unit_0.register_file_0.r13_10_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09890_ (
    .CLK(dco_clk),
    .D(_02008_),
    .Q(execution_unit_0.register_file_0.r13_11_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09891_ (
    .CLK(dco_clk),
    .D(_02009_),
    .Q(execution_unit_0.register_file_0.r13_12_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09892_ (
    .CLK(dco_clk),
    .D(_02010_),
    .Q(execution_unit_0.register_file_0.r13_13_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09893_ (
    .CLK(dco_clk),
    .D(_02011_),
    .Q(execution_unit_0.register_file_0.r13_14_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09894_ (
    .CLK(dco_clk),
    .D(_02012_),
    .Q(execution_unit_0.register_file_0.r13_15_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09895_ (
    .CLK(dco_clk),
    .D(_01990_),
    .Q(execution_unit_0.register_file_0.r12_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09896_ (
    .CLK(dco_clk),
    .D(_01997_),
    .Q(execution_unit_0.register_file_0.r12_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09897_ (
    .CLK(dco_clk),
    .D(_01998_),
    .Q(execution_unit_0.register_file_0.r12_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09898_ (
    .CLK(dco_clk),
    .D(_01999_),
    .Q(execution_unit_0.register_file_0.r12_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09899_ (
    .CLK(dco_clk),
    .D(_02000_),
    .Q(execution_unit_0.register_file_0.r12_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09900_ (
    .CLK(dco_clk),
    .D(_02001_),
    .Q(execution_unit_0.register_file_0.r12_5_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09901_ (
    .CLK(dco_clk),
    .D(_02002_),
    .Q(execution_unit_0.register_file_0.r12_6_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09902_ (
    .CLK(dco_clk),
    .D(_02003_),
    .Q(execution_unit_0.register_file_0.r12_7_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09903_ (
    .CLK(dco_clk),
    .D(_02004_),
    .Q(execution_unit_0.register_file_0.r12_8_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09904_ (
    .CLK(dco_clk),
    .D(_02005_),
    .Q(execution_unit_0.register_file_0.r12_9_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09905_ (
    .CLK(dco_clk),
    .D(_01991_),
    .Q(execution_unit_0.register_file_0.r12_10_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09906_ (
    .CLK(dco_clk),
    .D(_01992_),
    .Q(execution_unit_0.register_file_0.r12_11_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09907_ (
    .CLK(dco_clk),
    .D(_01993_),
    .Q(execution_unit_0.register_file_0.r12_12_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09908_ (
    .CLK(dco_clk),
    .D(_01994_),
    .Q(execution_unit_0.register_file_0.r12_13_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09909_ (
    .CLK(dco_clk),
    .D(_01995_),
    .Q(execution_unit_0.register_file_0.r12_14_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09910_ (
    .CLK(dco_clk),
    .D(_01996_),
    .Q(execution_unit_0.register_file_0.r12_15_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09911_ (
    .CLK(dco_clk),
    .D(_01974_),
    .Q(execution_unit_0.register_file_0.r11_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09912_ (
    .CLK(dco_clk),
    .D(_01981_),
    .Q(execution_unit_0.register_file_0.r11_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09913_ (
    .CLK(dco_clk),
    .D(_01982_),
    .Q(execution_unit_0.register_file_0.r11_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09914_ (
    .CLK(dco_clk),
    .D(_01983_),
    .Q(execution_unit_0.register_file_0.r11_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09915_ (
    .CLK(dco_clk),
    .D(_01984_),
    .Q(execution_unit_0.register_file_0.r11_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09916_ (
    .CLK(dco_clk),
    .D(_01985_),
    .Q(execution_unit_0.register_file_0.r11_5_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09917_ (
    .CLK(dco_clk),
    .D(_01986_),
    .Q(execution_unit_0.register_file_0.r11_6_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09918_ (
    .CLK(dco_clk),
    .D(_01987_),
    .Q(execution_unit_0.register_file_0.r11_7_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09919_ (
    .CLK(dco_clk),
    .D(_01988_),
    .Q(execution_unit_0.register_file_0.r11_8_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09920_ (
    .CLK(dco_clk),
    .D(_01989_),
    .Q(execution_unit_0.register_file_0.r11_9_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09921_ (
    .CLK(dco_clk),
    .D(_01975_),
    .Q(execution_unit_0.register_file_0.r11_10_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09922_ (
    .CLK(dco_clk),
    .D(_01976_),
    .Q(execution_unit_0.register_file_0.r11_11_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09923_ (
    .CLK(dco_clk),
    .D(_01977_),
    .Q(execution_unit_0.register_file_0.r11_12_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09924_ (
    .CLK(dco_clk),
    .D(_01978_),
    .Q(execution_unit_0.register_file_0.r11_13_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09925_ (
    .CLK(dco_clk),
    .D(_01979_),
    .Q(execution_unit_0.register_file_0.r11_14_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09926_ (
    .CLK(dco_clk),
    .D(_01980_),
    .Q(execution_unit_0.register_file_0.r11_15_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09927_ (
    .CLK(dco_clk),
    .D(_01958_),
    .Q(execution_unit_0.register_file_0.r10_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09928_ (
    .CLK(dco_clk),
    .D(_01965_),
    .Q(execution_unit_0.register_file_0.r10_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09929_ (
    .CLK(dco_clk),
    .D(_01966_),
    .Q(execution_unit_0.register_file_0.r10_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09930_ (
    .CLK(dco_clk),
    .D(_01967_),
    .Q(execution_unit_0.register_file_0.r10_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09931_ (
    .CLK(dco_clk),
    .D(_01968_),
    .Q(execution_unit_0.register_file_0.r10_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09932_ (
    .CLK(dco_clk),
    .D(_01969_),
    .Q(execution_unit_0.register_file_0.r10_5_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09933_ (
    .CLK(dco_clk),
    .D(_01970_),
    .Q(execution_unit_0.register_file_0.r10_6_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09934_ (
    .CLK(dco_clk),
    .D(_01971_),
    .Q(execution_unit_0.register_file_0.r10_7_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09935_ (
    .CLK(dco_clk),
    .D(_01972_),
    .Q(execution_unit_0.register_file_0.r10_8_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09936_ (
    .CLK(dco_clk),
    .D(_01973_),
    .Q(execution_unit_0.register_file_0.r10_9_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09937_ (
    .CLK(dco_clk),
    .D(_01959_),
    .Q(execution_unit_0.register_file_0.r10_10_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09938_ (
    .CLK(dco_clk),
    .D(_01960_),
    .Q(execution_unit_0.register_file_0.r10_11_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09939_ (
    .CLK(dco_clk),
    .D(_01961_),
    .Q(execution_unit_0.register_file_0.r10_12_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09940_ (
    .CLK(dco_clk),
    .D(_01962_),
    .Q(execution_unit_0.register_file_0.r10_13_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09941_ (
    .CLK(dco_clk),
    .D(_01963_),
    .Q(execution_unit_0.register_file_0.r10_14_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09942_ (
    .CLK(dco_clk),
    .D(_01964_),
    .Q(execution_unit_0.register_file_0.r10_15_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09943_ (
    .CLK(dco_clk),
    .D(_02174_),
    .Q(execution_unit_0.register_file_0.r9_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09944_ (
    .CLK(dco_clk),
    .D(_02181_),
    .Q(execution_unit_0.register_file_0.r9_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09945_ (
    .CLK(dco_clk),
    .D(_02182_),
    .Q(execution_unit_0.register_file_0.r9_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09946_ (
    .CLK(dco_clk),
    .D(_02183_),
    .Q(execution_unit_0.register_file_0.r9_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09947_ (
    .CLK(dco_clk),
    .D(_02184_),
    .Q(execution_unit_0.register_file_0.r9_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09948_ (
    .CLK(dco_clk),
    .D(_02185_),
    .Q(execution_unit_0.register_file_0.r9_5_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09949_ (
    .CLK(dco_clk),
    .D(_02186_),
    .Q(execution_unit_0.register_file_0.r9_6_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09950_ (
    .CLK(dco_clk),
    .D(_02187_),
    .Q(execution_unit_0.register_file_0.r9_7_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09951_ (
    .CLK(dco_clk),
    .D(_02188_),
    .Q(execution_unit_0.register_file_0.r9_8_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09952_ (
    .CLK(dco_clk),
    .D(_02189_),
    .Q(execution_unit_0.register_file_0.r9_9_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09953_ (
    .CLK(dco_clk),
    .D(_02175_),
    .Q(execution_unit_0.register_file_0.r9_10_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09954_ (
    .CLK(dco_clk),
    .D(_02176_),
    .Q(execution_unit_0.register_file_0.r9_11_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09955_ (
    .CLK(dco_clk),
    .D(_02177_),
    .Q(execution_unit_0.register_file_0.r9_12_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09956_ (
    .CLK(dco_clk),
    .D(_02178_),
    .Q(execution_unit_0.register_file_0.r9_13_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09957_ (
    .CLK(dco_clk),
    .D(_02179_),
    .Q(execution_unit_0.register_file_0.r9_14_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09958_ (
    .CLK(dco_clk),
    .D(_02180_),
    .Q(execution_unit_0.register_file_0.r9_15_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09959_ (
    .CLK(dco_clk),
    .D(_02158_),
    .Q(execution_unit_0.register_file_0.r8_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09960_ (
    .CLK(dco_clk),
    .D(_02165_),
    .Q(execution_unit_0.register_file_0.r8_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09961_ (
    .CLK(dco_clk),
    .D(_02166_),
    .Q(execution_unit_0.register_file_0.r8_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09962_ (
    .CLK(dco_clk),
    .D(_02167_),
    .Q(execution_unit_0.register_file_0.r8_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09963_ (
    .CLK(dco_clk),
    .D(_02168_),
    .Q(execution_unit_0.register_file_0.r8_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09964_ (
    .CLK(dco_clk),
    .D(_02169_),
    .Q(execution_unit_0.register_file_0.r8_5_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09965_ (
    .CLK(dco_clk),
    .D(_02170_),
    .Q(execution_unit_0.register_file_0.r8_6_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09966_ (
    .CLK(dco_clk),
    .D(_02171_),
    .Q(execution_unit_0.register_file_0.r8_7_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09967_ (
    .CLK(dco_clk),
    .D(_02172_),
    .Q(execution_unit_0.register_file_0.r8_8_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09968_ (
    .CLK(dco_clk),
    .D(_02173_),
    .Q(execution_unit_0.register_file_0.r8_9_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09969_ (
    .CLK(dco_clk),
    .D(_02159_),
    .Q(execution_unit_0.register_file_0.r8_10_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09970_ (
    .CLK(dco_clk),
    .D(_02160_),
    .Q(execution_unit_0.register_file_0.r8_11_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09971_ (
    .CLK(dco_clk),
    .D(_02161_),
    .Q(execution_unit_0.register_file_0.r8_12_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09972_ (
    .CLK(dco_clk),
    .D(_02162_),
    .Q(execution_unit_0.register_file_0.r8_13_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09973_ (
    .CLK(dco_clk),
    .D(_02163_),
    .Q(execution_unit_0.register_file_0.r8_14_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09974_ (
    .CLK(dco_clk),
    .D(_02164_),
    .Q(execution_unit_0.register_file_0.r8_15_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09975_ (
    .CLK(dco_clk),
    .D(_02142_),
    .Q(execution_unit_0.register_file_0.r7_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09976_ (
    .CLK(dco_clk),
    .D(_02149_),
    .Q(execution_unit_0.register_file_0.r7_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09977_ (
    .CLK(dco_clk),
    .D(_02150_),
    .Q(execution_unit_0.register_file_0.r7_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09978_ (
    .CLK(dco_clk),
    .D(_02151_),
    .Q(execution_unit_0.register_file_0.r7_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09979_ (
    .CLK(dco_clk),
    .D(_02152_),
    .Q(execution_unit_0.register_file_0.r7_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09980_ (
    .CLK(dco_clk),
    .D(_02153_),
    .Q(execution_unit_0.register_file_0.r7_5_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09981_ (
    .CLK(dco_clk),
    .D(_02154_),
    .Q(execution_unit_0.register_file_0.r7_6_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09982_ (
    .CLK(dco_clk),
    .D(_02155_),
    .Q(execution_unit_0.register_file_0.r7_7_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09983_ (
    .CLK(dco_clk),
    .D(_02156_),
    .Q(execution_unit_0.register_file_0.r7_8_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09984_ (
    .CLK(dco_clk),
    .D(_02157_),
    .Q(execution_unit_0.register_file_0.r7_9_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09985_ (
    .CLK(dco_clk),
    .D(_02143_),
    .Q(execution_unit_0.register_file_0.r7_10_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09986_ (
    .CLK(dco_clk),
    .D(_02144_),
    .Q(execution_unit_0.register_file_0.r7_11_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09987_ (
    .CLK(dco_clk),
    .D(_02145_),
    .Q(execution_unit_0.register_file_0.r7_12_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09988_ (
    .CLK(dco_clk),
    .D(_02146_),
    .Q(execution_unit_0.register_file_0.r7_13_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09989_ (
    .CLK(dco_clk),
    .D(_02147_),
    .Q(execution_unit_0.register_file_0.r7_14_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09990_ (
    .CLK(dco_clk),
    .D(_02148_),
    .Q(execution_unit_0.register_file_0.r7_15_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09991_ (
    .CLK(dco_clk),
    .D(_02126_),
    .Q(execution_unit_0.register_file_0.r6_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09992_ (
    .CLK(dco_clk),
    .D(_02133_),
    .Q(execution_unit_0.register_file_0.r6_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09993_ (
    .CLK(dco_clk),
    .D(_02134_),
    .Q(execution_unit_0.register_file_0.r6_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09994_ (
    .CLK(dco_clk),
    .D(_02135_),
    .Q(execution_unit_0.register_file_0.r6_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09995_ (
    .CLK(dco_clk),
    .D(_02136_),
    .Q(execution_unit_0.register_file_0.r6_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09996_ (
    .CLK(dco_clk),
    .D(_02137_),
    .Q(execution_unit_0.register_file_0.r6_5_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09997_ (
    .CLK(dco_clk),
    .D(_02138_),
    .Q(execution_unit_0.register_file_0.r6_6_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09998_ (
    .CLK(dco_clk),
    .D(_02139_),
    .Q(execution_unit_0.register_file_0.r6_7_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _09999_ (
    .CLK(dco_clk),
    .D(_02140_),
    .Q(execution_unit_0.register_file_0.r6_8_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10000_ (
    .CLK(dco_clk),
    .D(_02141_),
    .Q(execution_unit_0.register_file_0.r6_9_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10001_ (
    .CLK(dco_clk),
    .D(_02127_),
    .Q(execution_unit_0.register_file_0.r6_10_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10002_ (
    .CLK(dco_clk),
    .D(_02128_),
    .Q(execution_unit_0.register_file_0.r6_11_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10003_ (
    .CLK(dco_clk),
    .D(_02129_),
    .Q(execution_unit_0.register_file_0.r6_12_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10004_ (
    .CLK(dco_clk),
    .D(_02130_),
    .Q(execution_unit_0.register_file_0.r6_13_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10005_ (
    .CLK(dco_clk),
    .D(_02131_),
    .Q(execution_unit_0.register_file_0.r6_14_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10006_ (
    .CLK(dco_clk),
    .D(_02132_),
    .Q(execution_unit_0.register_file_0.r6_15_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10007_ (
    .CLK(dco_clk),
    .D(_02110_),
    .Q(execution_unit_0.register_file_0.r5_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10008_ (
    .CLK(dco_clk),
    .D(_02117_),
    .Q(execution_unit_0.register_file_0.r5_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10009_ (
    .CLK(dco_clk),
    .D(_02118_),
    .Q(execution_unit_0.register_file_0.r5_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10010_ (
    .CLK(dco_clk),
    .D(_02119_),
    .Q(execution_unit_0.register_file_0.r5_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10011_ (
    .CLK(dco_clk),
    .D(_02120_),
    .Q(execution_unit_0.register_file_0.r5_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10012_ (
    .CLK(dco_clk),
    .D(_02121_),
    .Q(execution_unit_0.register_file_0.r5_5_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10013_ (
    .CLK(dco_clk),
    .D(_02122_),
    .Q(execution_unit_0.register_file_0.r5_6_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10014_ (
    .CLK(dco_clk),
    .D(_02123_),
    .Q(execution_unit_0.register_file_0.r5_7_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10015_ (
    .CLK(dco_clk),
    .D(_02124_),
    .Q(execution_unit_0.register_file_0.r5_8_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10016_ (
    .CLK(dco_clk),
    .D(_02125_),
    .Q(execution_unit_0.register_file_0.r5_9_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10017_ (
    .CLK(dco_clk),
    .D(_02111_),
    .Q(execution_unit_0.register_file_0.r5_10_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10018_ (
    .CLK(dco_clk),
    .D(_02112_),
    .Q(execution_unit_0.register_file_0.r5_11_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10019_ (
    .CLK(dco_clk),
    .D(_02113_),
    .Q(execution_unit_0.register_file_0.r5_12_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10020_ (
    .CLK(dco_clk),
    .D(_02114_),
    .Q(execution_unit_0.register_file_0.r5_13_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10021_ (
    .CLK(dco_clk),
    .D(_02115_),
    .Q(execution_unit_0.register_file_0.r5_14_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10022_ (
    .CLK(dco_clk),
    .D(_02116_),
    .Q(execution_unit_0.register_file_0.r5_15_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10023_ (
    .CLK(dco_clk),
    .D(_02094_),
    .Q(execution_unit_0.register_file_0.r4_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10024_ (
    .CLK(dco_clk),
    .D(_02101_),
    .Q(execution_unit_0.register_file_0.r4_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10025_ (
    .CLK(dco_clk),
    .D(_02102_),
    .Q(execution_unit_0.register_file_0.r4_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10026_ (
    .CLK(dco_clk),
    .D(_02103_),
    .Q(execution_unit_0.register_file_0.r4_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10027_ (
    .CLK(dco_clk),
    .D(_02104_),
    .Q(execution_unit_0.register_file_0.r4_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10028_ (
    .CLK(dco_clk),
    .D(_02105_),
    .Q(execution_unit_0.register_file_0.r4_5_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10029_ (
    .CLK(dco_clk),
    .D(_02106_),
    .Q(execution_unit_0.register_file_0.r4_6_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10030_ (
    .CLK(dco_clk),
    .D(_02107_),
    .Q(execution_unit_0.register_file_0.r4_7_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10031_ (
    .CLK(dco_clk),
    .D(_02108_),
    .Q(execution_unit_0.register_file_0.r4_8_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10032_ (
    .CLK(dco_clk),
    .D(_02109_),
    .Q(execution_unit_0.register_file_0.r4_9_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10033_ (
    .CLK(dco_clk),
    .D(_02095_),
    .Q(execution_unit_0.register_file_0.r4_10_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10034_ (
    .CLK(dco_clk),
    .D(_02096_),
    .Q(execution_unit_0.register_file_0.r4_11_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10035_ (
    .CLK(dco_clk),
    .D(_02097_),
    .Q(execution_unit_0.register_file_0.r4_12_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10036_ (
    .CLK(dco_clk),
    .D(_02098_),
    .Q(execution_unit_0.register_file_0.r4_13_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10037_ (
    .CLK(dco_clk),
    .D(_02099_),
    .Q(execution_unit_0.register_file_0.r4_14_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10038_ (
    .CLK(dco_clk),
    .D(_02100_),
    .Q(execution_unit_0.register_file_0.r4_15_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10039_ (
    .CLK(dco_clk),
    .D(_02078_),
    .Q(execution_unit_0.register_file_0.r3_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10040_ (
    .CLK(dco_clk),
    .D(_02085_),
    .Q(execution_unit_0.register_file_0.r3_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10041_ (
    .CLK(dco_clk),
    .D(_02086_),
    .Q(execution_unit_0.register_file_0.r3_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10042_ (
    .CLK(dco_clk),
    .D(_02087_),
    .Q(execution_unit_0.register_file_0.r3_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10043_ (
    .CLK(dco_clk),
    .D(_02088_),
    .Q(execution_unit_0.register_file_0.r3_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10044_ (
    .CLK(dco_clk),
    .D(_02089_),
    .Q(execution_unit_0.register_file_0.r3_5_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10045_ (
    .CLK(dco_clk),
    .D(_02090_),
    .Q(execution_unit_0.register_file_0.r3_6_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10046_ (
    .CLK(dco_clk),
    .D(_02091_),
    .Q(execution_unit_0.register_file_0.r3_7_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10047_ (
    .CLK(dco_clk),
    .D(_02092_),
    .Q(execution_unit_0.register_file_0.r3_8_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10048_ (
    .CLK(dco_clk),
    .D(_02093_),
    .Q(execution_unit_0.register_file_0.r3_9_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10049_ (
    .CLK(dco_clk),
    .D(_02079_),
    .Q(execution_unit_0.register_file_0.r3_10_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10050_ (
    .CLK(dco_clk),
    .D(_02080_),
    .Q(execution_unit_0.register_file_0.r3_11_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10051_ (
    .CLK(dco_clk),
    .D(_02081_),
    .Q(execution_unit_0.register_file_0.r3_12_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10052_ (
    .CLK(dco_clk),
    .D(_02082_),
    .Q(execution_unit_0.register_file_0.r3_13_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10053_ (
    .CLK(dco_clk),
    .D(_02083_),
    .Q(execution_unit_0.register_file_0.r3_14_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10054_ (
    .CLK(dco_clk),
    .D(_02084_),
    .Q(execution_unit_0.register_file_0.r3_15_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10055_ (
    .CLK(dco_clk),
    .D(_02070_),
    .Q(execution_unit_0.alu_0.status_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10056_ (
    .CLK(dco_clk),
    .D(_02071_),
    .Q(execution_unit_0.alu_0.status_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10057_ (
    .CLK(dco_clk),
    .D(_02072_),
    .Q(execution_unit_0.alu_0.status_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10058_ (
    .CLK(dco_clk),
    .D(_02073_),
    .Q(execution_unit_0.gie ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10059_ (
    .CLK(dco_clk),
    .D(_02074_),
    .Q(execution_unit_0.register_file_0.r2_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10060_ (
    .CLK(dco_clk),
    .D(_02075_),
    .Q(clock_module_0.oscoff ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10061_ (
    .CLK(dco_clk),
    .D(_02076_),
    .Q(clock_module_0.scg1 ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10062_ (
    .CLK(dco_clk),
    .D(_02077_),
    .Q(execution_unit_0.alu_0.status_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10063_ (
    .CLK(dco_clk),
    .D(_02054_),
    .Q(execution_unit_0.register_file_0.r1_0_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10064_ (
    .CLK(dco_clk),
    .D(_02061_),
    .Q(execution_unit_0.register_file_0.r1_1_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10065_ (
    .CLK(dco_clk),
    .D(_02062_),
    .Q(execution_unit_0.register_file_0.r1_2_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10066_ (
    .CLK(dco_clk),
    .D(_02063_),
    .Q(execution_unit_0.register_file_0.r1_3_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10067_ (
    .CLK(dco_clk),
    .D(_02064_),
    .Q(execution_unit_0.register_file_0.r1_4_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10068_ (
    .CLK(dco_clk),
    .D(_02065_),
    .Q(execution_unit_0.register_file_0.r1_5_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10069_ (
    .CLK(dco_clk),
    .D(_02066_),
    .Q(execution_unit_0.register_file_0.r1_6_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10070_ (
    .CLK(dco_clk),
    .D(_02067_),
    .Q(execution_unit_0.register_file_0.r1_7_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10071_ (
    .CLK(dco_clk),
    .D(_02068_),
    .Q(execution_unit_0.register_file_0.r1_8_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10072_ (
    .CLK(dco_clk),
    .D(_02069_),
    .Q(execution_unit_0.register_file_0.r1_9_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10073_ (
    .CLK(dco_clk),
    .D(_02055_),
    .Q(execution_unit_0.register_file_0.r1_10_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10074_ (
    .CLK(dco_clk),
    .D(_02056_),
    .Q(execution_unit_0.register_file_0.r1_11_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10075_ (
    .CLK(dco_clk),
    .D(_02057_),
    .Q(execution_unit_0.register_file_0.r1_12_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10076_ (
    .CLK(dco_clk),
    .D(_02058_),
    .Q(execution_unit_0.register_file_0.r1_13_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10077_ (
    .CLK(dco_clk),
    .D(_02059_),
    .Q(execution_unit_0.register_file_0.r1_14_ ),
    .R(_02190_),
    .S(1'h1)
  );
  DFFSR _10078_ (
    .CLK(dco_clk),
    .D(_02060_),
    .Q(execution_unit_0.register_file_0.r1_15_ ),
    .R(_02190_),
    .S(1'h1)
  );
  INVX1 _10079_ (
    .A(e_state_3_),
    .Y(_03657_)
  );
  INVX1 _10080_ (
    .A(e_state_2_),
    .Y(_03658_)
  );
  INVX1 _10081_ (
    .A(e_state_0_),
    .Y(_03659_)
  );
  INVX1 _10082_ (
    .A(execution_unit_0.gie ),
    .Y(_03660_)
  );
  INVX1 _10083_ (
    .A(irq_13_),
    .Y(_03661_)
  );
  INVX1 _10084_ (
    .A(irq_7_),
    .Y(_03662_)
  );
  INVX1 _10085_ (
    .A(irq_3_),
    .Y(_03663_)
  );
  INVX1 _10086_ (
    .A(irq_1_),
    .Y(_03664_)
  );
  INVX1 _10087_ (
    .A(cpu_halt_cmd),
    .Y(_03665_)
  );
  INVX1 _10088_ (
    .A(1'h0),
    .Y(_03666_)
  );
  INVX1 _10089_ (
    .A(frontend_0.i_state_4_ ),
    .Y(_03667_)
  );
  INVX1 _10090_ (
    .A(frontend_0.exec_dst_wr ),
    .Y(_03668_)
  );
  INVX1 _10091_ (
    .A(frontend_0.exec_jmp ),
    .Y(_03669_)
  );
  INVX1 _10092_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .Y(_03670_)
  );
  INVX1 _10093_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .Y(_03671_)
  );
  INVX1 _10094_ (
    .A(dbg_0.fe_mdb_in_7_ ),
    .Y(_03672_)
  );
  INVX1 _10095_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .Y(_03673_)
  );
  INVX1 _10096_ (
    .A(dbg_0.fe_mdb_in_14_ ),
    .Y(_03674_)
  );
  INVX1 _10097_ (
    .A(dbg_0.fe_mdb_in_4_ ),
    .Y(_03675_)
  );
  INVX1 _10098_ (
    .A(dbg_0.fe_mdb_in_0_ ),
    .Y(_03676_)
  );
  INVX1 _10099_ (
    .A(dbg_0.fe_mdb_in_1_ ),
    .Y(_03677_)
  );
  INVX1 _10100_ (
    .A(dbg_0.fe_mdb_in_2_ ),
    .Y(_03678_)
  );
  INVX1 _10101_ (
    .A(dbg_0.fe_mdb_in_3_ ),
    .Y(_03679_)
  );
  INVX1 _10102_ (
    .A(execution_unit_0.UNUSED_inst_ad_idx ),
    .Y(_03680_)
  );
  INVX1 _10103_ (
    .A(frontend_0.i_state_5_ ),
    .Y(_03681_)
  );
  INVX1 _10104_ (
    .A(frontend_0.i_state_2_ ),
    .Y(_03682_)
  );
  INVX1 _10105_ (
    .A(execution_unit_0.pc_sw_wr ),
    .Y(_03683_)
  );
  INVX1 _10106_ (
    .A(frontend_0.inst_sz_0_ ),
    .Y(_03684_)
  );
  INVX1 _10107_ (
    .A(frontend_0.i_state_1_ ),
    .Y(_03685_)
  );
  INVX1 _10108_ (
    .A(frontend_0.i_state_3_ ),
    .Y(_03686_)
  );
  INVX1 _10109_ (
    .A(frontend_0.i_state_0_ ),
    .Y(_03687_)
  );
  INVX1 _10110_ (
    .A(execution_unit_0.alu_0.alu_out_0_ ),
    .Y(_03688_)
  );
  INVX1 _10111_ (
    .A(dbg_0.UNUSED_pc_1_ ),
    .Y(_03689_)
  );
  INVX1 _10112_ (
    .A(frontend_0.irq_addr_1_ ),
    .Y(_03690_)
  );
  INVX1 _10113_ (
    .A(dbg_0.UNUSED_pc_2_ ),
    .Y(_03691_)
  );
  INVX1 _10114_ (
    .A(frontend_0.irq_addr_2_ ),
    .Y(_03692_)
  );
  INVX1 _10115_ (
    .A(dbg_0.UNUSED_pc_3_ ),
    .Y(_03693_)
  );
  INVX1 _10116_ (
    .A(frontend_0.irq_addr_3_ ),
    .Y(_03694_)
  );
  INVX1 _10117_ (
    .A(dbg_0.UNUSED_pc_4_ ),
    .Y(_03695_)
  );
  INVX1 _10118_ (
    .A(dbg_0.UNUSED_pc_5_ ),
    .Y(_03696_)
  );
  INVX1 _10119_ (
    .A(dbg_0.UNUSED_pc_6_ ),
    .Y(_03697_)
  );
  INVX1 _10120_ (
    .A(dbg_0.fe_mdb_in_6_ ),
    .Y(_03698_)
  );
  INVX1 _10121_ (
    .A(frontend_0.irq_addr_6_ ),
    .Y(_03699_)
  );
  INVX1 _10122_ (
    .A(dbg_0.UNUSED_pc_7_ ),
    .Y(_03700_)
  );
  INVX1 _10123_ (
    .A(dbg_0.UNUSED_pc_8_ ),
    .Y(_03701_)
  );
  INVX1 _10124_ (
    .A(dbg_0.UNUSED_pc_9_ ),
    .Y(_03702_)
  );
  INVX1 _10125_ (
    .A(dbg_0.UNUSED_pc_10_ ),
    .Y(_03703_)
  );
  INVX1 _10126_ (
    .A(dbg_0.UNUSED_pc_11_ ),
    .Y(_03704_)
  );
  INVX1 _10127_ (
    .A(dbg_0.UNUSED_pc_12_ ),
    .Y(_03705_)
  );
  INVX1 _10128_ (
    .A(dbg_0.fe_mdb_in_12_ ),
    .Y(_03706_)
  );
  INVX1 _10129_ (
    .A(dbg_0.UNUSED_pc_13_ ),
    .Y(_03707_)
  );
  INVX1 _10130_ (
    .A(dbg_0.UNUSED_pc_14_ ),
    .Y(_03708_)
  );
  INVX1 _10131_ (
    .A(dbg_0.UNUSED_pc_15_ ),
    .Y(_03709_)
  );
  INVX1 _10132_ (
    .A(frontend_0.inst_dest_bin_3_ ),
    .Y(_03710_)
  );
  INVX1 _10133_ (
    .A(frontend_0.inst_dest_bin_2_ ),
    .Y(_03711_)
  );
  INVX1 _10134_ (
    .A(frontend_0.inst_dest_bin_0_ ),
    .Y(_03712_)
  );
  INVX1 _10135_ (
    .A(frontend_0.inst_dest_bin_1_ ),
    .Y(_03713_)
  );
  INVX1 _10136_ (
    .A(execution_unit_0.inst_type_1_ ),
    .Y(_03714_)
  );
  INVX1 _10137_ (
    .A(dbg_0.dbg_mem_addr_0_ ),
    .Y(_03715_)
  );
  INVX1 _10138_ (
    .A(dbg_0.dbg_mem_addr_1_ ),
    .Y(_03716_)
  );
  INVX1 _10139_ (
    .A(dbg_0.dbg_mem_addr_3_ ),
    .Y(_03717_)
  );
  INVX1 _10140_ (
    .A(dbg_0.dbg_mem_addr_2_ ),
    .Y(_03718_)
  );
  INVX1 _10141_ (
    .A(execution_unit_0.inst_type_0_ ),
    .Y(_03719_)
  );
  INVX1 _10142_ (
    .A(frontend_0.inst_src_bin_1_ ),
    .Y(_03720_)
  );
  INVX1 _10143_ (
    .A(frontend_0.inst_src_bin_3_ ),
    .Y(_03721_)
  );
  INVX1 _10144_ (
    .A(frontend_0.inst_src_bin_2_ ),
    .Y(_03722_)
  );
  INVX1 _10145_ (
    .A(execution_unit_0.inst_type_2_ ),
    .Y(_03723_)
  );
  INVX1 _10146_ (
    .A(execution_unit_0.alu_0.inst_alu_3_ ),
    .Y(_03724_)
  );
  INVX1 _10147_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_03725_)
  );
  INVX1 _10148_ (
    .A(execution_unit_0.alu_0.inst_alu_8_ ),
    .Y(_03726_)
  );
  INVX1 _10149_ (
    .A(frontend_0.inst_jmp_bin_0_ ),
    .Y(_03727_)
  );
  INVX1 _10150_ (
    .A(frontend_0.inst_jmp_bin_1_ ),
    .Y(_03728_)
  );
  INVX1 _10151_ (
    .A(execution_unit_0.inst_irq_rst ),
    .Y(_03729_)
  );
  INVX1 _10152_ (
    .A(_00162_),
    .Y(_03438_)
  );
  NOR2X1 _10153_ (
    .A(e_state_0_),
    .B(e_state_1_),
    .Y(_03730_)
  );
  INVX1 _10154_ (
    .A(_03730_),
    .Y(_03731_)
  );
  NAND2X1 _10155_ (
    .A(e_state_3_),
    .B(e_state_2_),
    .Y(_03732_)
  );
  OAI21X1 _10156_ (
    .A(_03731_),
    .B(_03732_),
    .C(frontend_0.exec_jmp ),
    .Y(_03733_)
  );
  INVX1 _10157_ (
    .A(_03733_),
    .Y(_03734_)
  );
  NOR2X1 _10158_ (
    .A(_03657_),
    .B(e_state_2_),
    .Y(_03735_)
  );
  NAND2X1 _10159_ (
    .A(e_state_3_),
    .B(_03658_),
    .Y(_03736_)
  );
  NAND2X1 _10160_ (
    .A(_03659_),
    .B(e_state_1_),
    .Y(_03737_)
  );
  NOR2X1 _10161_ (
    .A(_03736_),
    .B(_03737_),
    .Y(_03738_)
  );
  OR2X1 _10162_ (
    .A(_03736_),
    .B(_03737_),
    .Y(_03739_)
  );
  OAI21X1 _10163_ (
    .A(_03736_),
    .B(_03737_),
    .C(frontend_0.exec_dst_wr ),
    .Y(_03740_)
  );
  AND2X1 _10164_ (
    .A(e_state_0_),
    .B(e_state_1_),
    .Y(_03741_)
  );
  NAND2X1 _10165_ (
    .A(e_state_0_),
    .B(e_state_1_),
    .Y(_03742_)
  );
  NAND2X1 _10166_ (
    .A(_03657_),
    .B(e_state_2_),
    .Y(_03743_)
  );
  NOR2X1 _10167_ (
    .A(_03742_),
    .B(_03743_),
    .Y(_03744_)
  );
  NAND3X1 _10168_ (
    .A(_03657_),
    .B(e_state_2_),
    .C(_03741_),
    .Y(_03745_)
  );
  NAND3X1 _10169_ (
    .A(e_state_3_),
    .B(_03658_),
    .C(_03741_),
    .Y(_03746_)
  );
  MUX2X1 _10170_ (
    .A(_03745_),
    .B(_03746_),
    .S(frontend_0.exec_src_wr ),
    .Y(_03747_)
  );
  OAI21X1 _10171_ (
    .A(frontend_0.exec_dst_wr ),
    .B(_03747_),
    .C(_03740_),
    .Y(_03748_)
  );
  AOI21X1 _10172_ (
    .A(_03669_),
    .B(_03748_),
    .C(_03734_),
    .Y(exec_done)
  );
  NOR2X1 _10173_ (
    .A(frontend_0.i_state_4_ ),
    .B(exec_done),
    .Y(_03749_)
  );
  NOR2X1 _10174_ (
    .A(irq_12_),
    .B(irq_13_),
    .Y(_03750_)
  );
  NOR2X1 _10175_ (
    .A(irq_6_),
    .B(irq_7_),
    .Y(_03751_)
  );
  NOR2X1 _10176_ (
    .A(frontend_0.wdt_irq ),
    .B(irq_10_),
    .Y(_03752_)
  );
  NOR2X1 _10177_ (
    .A(irq_11_),
    .B(irq_9_),
    .Y(_03753_)
  );
  NAND2X1 _10178_ (
    .A(_03752_),
    .B(_03753_),
    .Y(_03754_)
  );
  NOR2X1 _10179_ (
    .A(irq_8_),
    .B(irq_2_),
    .Y(_03755_)
  );
  NAND3X1 _10180_ (
    .A(_03663_),
    .B(_03664_),
    .C(_03755_),
    .Y(_03756_)
  );
  NOR3X1 _10181_ (
    .A(irq_4_),
    .B(irq_5_),
    .C(irq_0_),
    .Y(_03757_)
  );
  NAND3X1 _10182_ (
    .A(_03750_),
    .B(_03751_),
    .C(_03757_),
    .Y(_03758_)
  );
  NOR3X1 _10183_ (
    .A(_03754_),
    .B(_03756_),
    .C(_03758_),
    .Y(_03759_)
  );
  OAI21X1 _10184_ (
    .A(_03660_),
    .B(_03759_),
    .C(_03666_),
    .Y(_03760_)
  );
  AND2X1 _10185_ (
    .A(cpu_en),
    .B(_03665_),
    .Y(_03761_)
  );
  NAND2X1 _10186_ (
    .A(cpu_en),
    .B(_03665_),
    .Y(_03762_)
  );
  NOR2X1 _10187_ (
    .A(cpu_halt_st),
    .B(_03762_),
    .Y(_03763_)
  );
  AND2X1 _10188_ (
    .A(_03760_),
    .B(_03763_),
    .Y(_03764_)
  );
  NAND2X1 _10189_ (
    .A(_03760_),
    .B(_03763_),
    .Y(_03765_)
  );
  NOR2X1 _10190_ (
    .A(_03749_),
    .B(_03765_),
    .Y(_03766_)
  );
  OAI21X1 _10191_ (
    .A(frontend_0.i_state_4_ ),
    .B(exec_done),
    .C(_03764_),
    .Y(_03767_)
  );
  NOR2X1 _10192_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(dbg_0.fe_mdb_in_14_ ),
    .Y(_03768_)
  );
  OAI21X1 _10193_ (
    .A(_03749_),
    .B(_03765_),
    .C(_03768_),
    .Y(_03769_)
  );
  NOR2X1 _10194_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(_03769_),
    .Y(_03770_)
  );
  NAND3X1 _10195_ (
    .A(_03673_),
    .B(_03767_),
    .C(_03768_),
    .Y(_03771_)
  );
  NAND2X1 _10196_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(dbg_0.fe_mdb_in_7_ ),
    .Y(_03772_)
  );
  NOR2X1 _10197_ (
    .A(_03771_),
    .B(_03772_),
    .Y(_03773_)
  );
  OR2X1 _10198_ (
    .A(_03771_),
    .B(_03772_),
    .Y(_03774_)
  );
  AOI21X1 _10199_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(_03773_),
    .C(_03766_),
    .Y(_03775_)
  );
  NOR2X1 _10200_ (
    .A(cpu_halt_st),
    .B(_03775_),
    .Y(_03776_)
  );
  OR2X1 _10201_ (
    .A(cpu_halt_st),
    .B(_03775_),
    .Y(_03777_)
  );
  OR2X1 _10202_ (
    .A(_03673_),
    .B(_03769_),
    .Y(_03778_)
  );
  INVX1 _10203_ (
    .A(_03778_),
    .Y(_03779_)
  );
  AND2X1 _10204_ (
    .A(dbg_0.fe_mdb_in_5_ ),
    .B(_03778_),
    .Y(_03780_)
  );
  OAI21X1 _10205_ (
    .A(_03673_),
    .B(_03769_),
    .C(dbg_0.fe_mdb_in_5_ ),
    .Y(_03781_)
  );
  NAND2X1 _10206_ (
    .A(dbg_0.fe_mdb_in_4_ ),
    .B(_03780_),
    .Y(_03782_)
  );
  NOR2X1 _10207_ (
    .A(dbg_0.fe_mdb_in_2_ ),
    .B(dbg_0.fe_mdb_in_3_ ),
    .Y(_03783_)
  );
  NAND2X1 _10208_ (
    .A(_03678_),
    .B(_03679_),
    .Y(_03784_)
  );
  NOR2X1 _10209_ (
    .A(dbg_0.fe_mdb_in_10_ ),
    .B(dbg_0.fe_mdb_in_11_ ),
    .Y(_03785_)
  );
  INVX1 _10210_ (
    .A(_03785_),
    .Y(_03786_)
  );
  MUX2X1 _10211_ (
    .A(_03786_),
    .B(_03784_),
    .S(_03771_),
    .Y(_03787_)
  );
  MUX2X1 _10212_ (
    .A(_03785_),
    .B(_03783_),
    .S(_03771_),
    .Y(_03788_)
  );
  MUX2X1 _10213_ (
    .A(_03670_),
    .B(_03677_),
    .S(_03771_),
    .Y(_03789_)
  );
  MUX2X1 _10214_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(dbg_0.fe_mdb_in_1_ ),
    .S(_03771_),
    .Y(_03790_)
  );
  NOR2X1 _10215_ (
    .A(_03788_),
    .B(_03790_),
    .Y(_03791_)
  );
  NAND2X1 _10216_ (
    .A(_03787_),
    .B(_03789_),
    .Y(_03792_)
  );
  NOR2X1 _10217_ (
    .A(_03782_),
    .B(_03791_),
    .Y(_03793_)
  );
  NAND2X1 _10218_ (
    .A(_03675_),
    .B(_03780_),
    .Y(_03794_)
  );
  NAND2X1 _10219_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(_03672_),
    .Y(_03795_)
  );
  NOR2X1 _10220_ (
    .A(_03771_),
    .B(_03795_),
    .Y(_03796_)
  );
  INVX1 _10221_ (
    .A(_03796_),
    .Y(_03797_)
  );
  NAND2X1 _10222_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(_03796_),
    .Y(_03798_)
  );
  MUX2X1 _10223_ (
    .A(_03671_),
    .B(_03676_),
    .S(_03771_),
    .Y(_03799_)
  );
  MUX2X1 _10224_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(dbg_0.fe_mdb_in_0_ ),
    .S(_03771_),
    .Y(_03800_)
  );
  NAND3X1 _10225_ (
    .A(_03787_),
    .B(_03790_),
    .C(_03800_),
    .Y(_03801_)
  );
  NAND2X1 _10226_ (
    .A(_03793_),
    .B(_03801_),
    .Y(_03802_)
  );
  OR2X1 _10227_ (
    .A(_03782_),
    .B(_03801_),
    .Y(_03803_)
  );
  AOI22X1 _10228_ (
    .A(_03780_),
    .B(_03792_),
    .C(_03796_),
    .D(dbg_0.fe_mdb_in_8_ ),
    .Y(_03804_)
  );
  OAI21X1 _10229_ (
    .A(_03781_),
    .B(_03791_),
    .C(_03798_),
    .Y(_03805_)
  );
  NOR2X1 _10230_ (
    .A(_03766_),
    .B(_03768_),
    .Y(_03806_)
  );
  NAND2X1 _10231_ (
    .A(dbg_0.fe_mdb_in_7_ ),
    .B(_03806_),
    .Y(_03807_)
  );
  NOR2X1 _10232_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(_03771_),
    .Y(_03808_)
  );
  NAND2X1 _10233_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(_03808_),
    .Y(_03809_)
  );
  AOI21X1 _10234_ (
    .A(_03807_),
    .B(_03809_),
    .C(_03805_),
    .Y(_03810_)
  );
  OR2X1 _10235_ (
    .A(clock_module_0.UNUSED_cpuoff ),
    .B(_03762_),
    .Y(_03811_)
  );
  NOR2X1 _10236_ (
    .A(frontend_0.i_state_4_ ),
    .B(_03811_),
    .Y(_03812_)
  );
  OR2X1 _10237_ (
    .A(frontend_0.i_state_4_ ),
    .B(_03811_),
    .Y(_03813_)
  );
  NOR3X1 _10238_ (
    .A(_03788_),
    .B(_03790_),
    .C(_03800_),
    .Y(_03814_)
  );
  NAND3X1 _10239_ (
    .A(_03787_),
    .B(_03789_),
    .C(_03799_),
    .Y(_03815_)
  );
  OAI21X1 _10240_ (
    .A(_03673_),
    .B(_03769_),
    .C(dbg_0.fe_mdb_in_4_ ),
    .Y(_03816_)
  );
  NOR2X1 _10241_ (
    .A(dbg_0.fe_mdb_in_5_ ),
    .B(_03816_),
    .Y(_03817_)
  );
  OR2X1 _10242_ (
    .A(dbg_0.fe_mdb_in_5_ ),
    .B(_03816_),
    .Y(_03818_)
  );
  OAI21X1 _10243_ (
    .A(_03792_),
    .B(_03800_),
    .C(_03817_),
    .Y(_03819_)
  );
  AOI21X1 _10244_ (
    .A(_03815_),
    .B(_03817_),
    .C(_03813_),
    .Y(_03820_)
  );
  OAI21X1 _10245_ (
    .A(_03814_),
    .B(_03818_),
    .C(_03812_),
    .Y(_03821_)
  );
  OAI21X1 _10246_ (
    .A(_03810_),
    .B(_03821_),
    .C(_03777_),
    .Y(_03822_)
  );
  NOR2X1 _10247_ (
    .A(frontend_0.exec_jmp ),
    .B(_03746_),
    .Y(_03823_)
  );
  NOR2X1 _10248_ (
    .A(e_state_1_),
    .B(_03732_),
    .Y(_03824_)
  );
  NOR2X1 _10249_ (
    .A(_03744_),
    .B(_03824_),
    .Y(_03825_)
  );
  OAI21X1 _10250_ (
    .A(frontend_0.exec_jmp ),
    .B(_03739_),
    .C(_03825_),
    .Y(_03826_)
  );
  OAI21X1 _10251_ (
    .A(_03823_),
    .B(_03826_),
    .C(_03822_),
    .Y(_03827_)
  );
  OR2X1 _10252_ (
    .A(_03659_),
    .B(e_state_1_),
    .Y(_03828_)
  );
  NOR2X1 _10253_ (
    .A(_03736_),
    .B(_03828_),
    .Y(_03829_)
  );
  NOR2X1 _10254_ (
    .A(_03731_),
    .B(_03743_),
    .Y(_03830_)
  );
  NOR2X1 _10255_ (
    .A(_03829_),
    .B(_03830_),
    .Y(_03831_)
  );
  OAI21X1 _10256_ (
    .A(_03668_),
    .B(_03746_),
    .C(_03831_),
    .Y(_03832_)
  );
  NAND2X1 _10257_ (
    .A(_03657_),
    .B(_03658_),
    .Y(_03833_)
  );
  OR2X1 _10258_ (
    .A(e_state_0_),
    .B(_03833_),
    .Y(_03834_)
  );
  MUX2X1 _10259_ (
    .A(_03732_),
    .B(_03834_),
    .S(e_state_1_),
    .Y(_03835_)
  );
  NOR2X1 _10260_ (
    .A(_03832_),
    .B(_03835_),
    .Y(_03836_)
  );
  NOR2X1 _10261_ (
    .A(_03737_),
    .B(_03743_),
    .Y(_03837_)
  );
  NOR2X1 _10262_ (
    .A(execution_unit_0.UNUSED_inst_ad_symb ),
    .B(execution_unit_0.inst_ad_6_ ),
    .Y(_03838_)
  );
  NAND3X1 _10263_ (
    .A(_03680_),
    .B(_03837_),
    .C(_03838_),
    .Y(_03839_)
  );
  OR2X1 _10264_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .B(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .Y(_03840_)
  );
  OR2X1 _10265_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_03840_),
    .Y(_03841_)
  );
  NAND2X1 _10266_ (
    .A(frontend_0.exec_src_wr ),
    .B(_03823_),
    .Y(_03842_)
  );
  OAI21X1 _10267_ (
    .A(_03839_),
    .B(_03841_),
    .C(_03842_),
    .Y(_03843_)
  );
  NOR2X1 _10268_ (
    .A(execution_unit_0.inst_as_4_ ),
    .B(execution_unit_0.inst_as_1_ ),
    .Y(_03844_)
  );
  NOR2X1 _10269_ (
    .A(execution_unit_0.inst_as_6_ ),
    .B(execution_unit_0.inst_as_5_ ),
    .Y(_03845_)
  );
  NAND2X1 _10270_ (
    .A(_03844_),
    .B(_03845_),
    .Y(_03846_)
  );
  INVX1 _10271_ (
    .A(_03846_),
    .Y(_03847_)
  );
  NOR2X1 _10272_ (
    .A(_03681_),
    .B(_03847_),
    .Y(_03848_)
  );
  INVX1 _10273_ (
    .A(_03848_),
    .Y(_03849_)
  );
  OR2X1 _10274_ (
    .A(_03743_),
    .B(_03828_),
    .Y(_03850_)
  );
  INVX1 _10275_ (
    .A(_03850_),
    .Y(_03851_)
  );
  AOI21X1 _10276_ (
    .A(_03848_),
    .B(_03851_),
    .C(_03843_),
    .Y(_03852_)
  );
  NAND3X1 _10277_ (
    .A(_03827_),
    .B(_03836_),
    .C(_03852_),
    .Y(frontend_0.e_state_nxt_1_ )
  );
  OAI21X1 _10278_ (
    .A(frontend_0.i_state_4_ ),
    .B(frontend_0.i_state_2_ ),
    .C(_03766_),
    .Y(_03853_)
  );
  INVX1 _10279_ (
    .A(_03853_),
    .Y(_03434_)
  );
  NAND2X1 _10280_ (
    .A(e_state_0_),
    .B(_03824_),
    .Y(_03854_)
  );
  NOR2X1 _10281_ (
    .A(_03761_),
    .B(_03854_),
    .Y(_03855_)
  );
  OAI21X1 _10282_ (
    .A(exec_done),
    .B(_03855_),
    .C(_03811_),
    .Y(_03856_)
  );
  NAND3X1 _10283_ (
    .A(frontend_0.i_state_2_ ),
    .B(_03767_),
    .C(_03856_),
    .Y(_03857_)
  );
  AOI21X1 _10284_ (
    .A(_03681_),
    .B(_03857_),
    .C(_03683_),
    .Y(_03858_)
  );
  NAND3X1 _10285_ (
    .A(_03683_),
    .B(_03767_),
    .C(_03856_),
    .Y(_03859_)
  );
  INVX1 _10286_ (
    .A(_03859_),
    .Y(_03860_)
  );
  AOI21X1 _10287_ (
    .A(e_state_0_),
    .B(_03824_),
    .C(exec_done),
    .Y(_03861_)
  );
  NAND2X1 _10288_ (
    .A(frontend_0.i_state_2_ ),
    .B(_03861_),
    .Y(_03862_)
  );
  INVX1 _10289_ (
    .A(_03862_),
    .Y(_03863_)
  );
  NOR2X1 _10290_ (
    .A(_03667_),
    .B(_03811_),
    .Y(_03864_)
  );
  OR2X1 _10291_ (
    .A(_03684_),
    .B(frontend_0.inst_sz_1_ ),
    .Y(_03865_)
  );
  NOR2X1 _10292_ (
    .A(_03681_),
    .B(execution_unit_0.pc_sw_wr ),
    .Y(_03866_)
  );
  INVX1 _10293_ (
    .A(_03866_),
    .Y(_03867_)
  );
  NOR2X1 _10294_ (
    .A(frontend_0.i_state_1_ ),
    .B(frontend_0.i_state_3_ ),
    .Y(_03868_)
  );
  OAI21X1 _10295_ (
    .A(_03865_),
    .B(_03867_),
    .C(_03868_),
    .Y(_03869_)
  );
  AOI21X1 _10296_ (
    .A(_03765_),
    .B(_03864_),
    .C(_03869_),
    .Y(_03870_)
  );
  OAI21X1 _10297_ (
    .A(_03859_),
    .B(_03862_),
    .C(_03870_),
    .Y(_03871_)
  );
  NOR2X1 _10298_ (
    .A(_03858_),
    .B(_03871_),
    .Y(_03872_)
  );
  NOR2X1 _10299_ (
    .A(_03682_),
    .B(_03861_),
    .Y(dbg_0.decode_noirq )
  );
  NAND2X1 _10300_ (
    .A(_03860_),
    .B(dbg_0.decode_noirq ),
    .Y(_03873_)
  );
  NAND2X1 _10301_ (
    .A(_03872_),
    .B(_03873_),
    .Y(_03874_)
  );
  AND2X1 _10302_ (
    .A(_03803_),
    .B(_03819_),
    .Y(_03875_)
  );
  AND2X1 _10303_ (
    .A(_03807_),
    .B(_03875_),
    .Y(_03876_)
  );
  INVX1 _10304_ (
    .A(_03876_),
    .Y(_03877_)
  );
  OAI21X1 _10305_ (
    .A(_03873_),
    .B(_03877_),
    .C(_03872_),
    .Y(_03435_)
  );
  NAND2X1 _10306_ (
    .A(frontend_0.i_state_2_ ),
    .B(_03855_),
    .Y(_03878_)
  );
  OAI21X1 _10307_ (
    .A(frontend_0.i_state_4_ ),
    .B(frontend_0.i_state_2_ ),
    .C(_03811_),
    .Y(_03879_)
  );
  OR2X1 _10308_ (
    .A(_03764_),
    .B(_03879_),
    .Y(_03880_)
  );
  OAI21X1 _10309_ (
    .A(_03749_),
    .B(_03880_),
    .C(_03878_),
    .Y(_03436_)
  );
  NOR2X1 _10310_ (
    .A(_03873_),
    .B(_03876_),
    .Y(_03433_)
  );
  OAI21X1 _10311_ (
    .A(_03684_),
    .B(frontend_0.inst_sz_1_ ),
    .C(_03866_),
    .Y(_03881_)
  );
  INVX1 _10312_ (
    .A(_03881_),
    .Y(_03432_)
  );
  NAND2X1 _10313_ (
    .A(_03683_),
    .B(_03687_),
    .Y(_03882_)
  );
  AOI21X1 _10314_ (
    .A(_03676_),
    .B(frontend_0.i_state_3_ ),
    .C(_03882_),
    .Y(_03883_)
  );
  OAI21X1 _10315_ (
    .A(frontend_0.i_state_3_ ),
    .B(dbg_0.UNUSED_pc_0_ ),
    .C(_03883_),
    .Y(_03884_)
  );
  OAI21X1 _10316_ (
    .A(_03683_),
    .B(_03688_),
    .C(_03884_),
    .Y(UNUSED_fe_mab_0)
  );
  AOI21X1 _10317_ (
    .A(_03804_),
    .B(_03820_),
    .C(_03776_),
    .Y(_03885_)
  );
  OAI21X1 _10318_ (
    .A(_03805_),
    .B(_03821_),
    .C(_03777_),
    .Y(_03886_)
  );
  NOR3X1 _10319_ (
    .A(frontend_0.exec_src_wr ),
    .B(frontend_0.exec_jmp ),
    .C(_03885_),
    .Y(_03887_)
  );
  NOR2X1 _10320_ (
    .A(frontend_0.exec_dst_wr ),
    .B(_03746_),
    .Y(_03888_)
  );
  INVX1 _10321_ (
    .A(_03888_),
    .Y(_03889_)
  );
  NOR2X1 _10322_ (
    .A(_03887_),
    .B(_03889_),
    .Y(_03890_)
  );
  OR2X1 _10323_ (
    .A(_03887_),
    .B(_03889_),
    .Y(_03891_)
  );
  AOI21X1 _10324_ (
    .A(_03669_),
    .B(_03886_),
    .C(_03739_),
    .Y(_03892_)
  );
  NOR2X1 _10325_ (
    .A(_03742_),
    .B(_03833_),
    .Y(_03893_)
  );
  NOR2X1 _10326_ (
    .A(_03851_),
    .B(_03893_),
    .Y(_03894_)
  );
  OAI21X1 _10327_ (
    .A(_03825_),
    .B(_03886_),
    .C(_03894_),
    .Y(_03895_)
  );
  NOR2X1 _10328_ (
    .A(_03892_),
    .B(_03895_),
    .Y(_03896_)
  );
  OR2X1 _10329_ (
    .A(_03892_),
    .B(_03895_),
    .Y(_03897_)
  );
  OAI21X1 _10330_ (
    .A(_03887_),
    .B(_03889_),
    .C(_03896_),
    .Y(frontend_0.e_state_nxt_2_ )
  );
  NOR2X1 _10331_ (
    .A(_03683_),
    .B(execution_unit_0.alu_0.alu_out_1_ ),
    .Y(_03898_)
  );
  AOI21X1 _10332_ (
    .A(_03804_),
    .B(_03819_),
    .C(_03813_),
    .Y(_03899_)
  );
  OAI21X1 _10333_ (
    .A(frontend_0.exec_src_wr ),
    .B(_03746_),
    .C(_03825_),
    .Y(_03900_)
  );
  OAI21X1 _10334_ (
    .A(_03738_),
    .B(_03900_),
    .C(_03777_),
    .Y(_03901_)
  );
  NAND2X1 _10335_ (
    .A(e_state_1_),
    .B(frontend_0.exec_jmp ),
    .Y(_03902_)
  );
  NAND2X1 _10336_ (
    .A(_03730_),
    .B(_03735_),
    .Y(_03903_)
  );
  AOI21X1 _10337_ (
    .A(_03730_),
    .B(_03735_),
    .C(_03837_),
    .Y(_03904_)
  );
  OAI21X1 _10338_ (
    .A(_03736_),
    .B(_03902_),
    .C(_03904_),
    .Y(_03905_)
  );
  NOR2X1 _10339_ (
    .A(_03832_),
    .B(_03905_),
    .Y(_03906_)
  );
  OAI21X1 _10340_ (
    .A(_03899_),
    .B(_03901_),
    .C(_03906_),
    .Y(frontend_0.e_state_nxt_3_ )
  );
  AOI21X1 _10341_ (
    .A(_03804_),
    .B(_03807_),
    .C(_03821_),
    .Y(_03907_)
  );
  AND2X1 _10342_ (
    .A(_03668_),
    .B(_03823_),
    .Y(_03908_)
  );
  OAI21X1 _10343_ (
    .A(_03826_),
    .B(_03908_),
    .C(_03777_),
    .Y(_03909_)
  );
  AOI21X1 _10344_ (
    .A(frontend_0.i_state_5_ ),
    .B(_03847_),
    .C(frontend_0.i_state_1_ ),
    .Y(_03910_)
  );
  INVX1 _10345_ (
    .A(_03910_),
    .Y(_03911_)
  );
  NOR2X1 _10346_ (
    .A(frontend_0.exec_dext_rdy ),
    .B(_03911_),
    .Y(_03912_)
  );
  NOR2X1 _10347_ (
    .A(_03903_),
    .B(_03912_),
    .Y(_03913_)
  );
  NAND3X1 _10348_ (
    .A(_03831_),
    .B(_03834_),
    .C(_03839_),
    .Y(_03914_)
  );
  AOI21X1 _10349_ (
    .A(_03849_),
    .B(_03851_),
    .C(_03914_),
    .Y(_03915_)
  );
  OAI21X1 _10350_ (
    .A(frontend_0.exec_dst_wr ),
    .B(_03842_),
    .C(_03915_),
    .Y(_03916_)
  );
  NOR2X1 _10351_ (
    .A(_03913_),
    .B(_03916_),
    .Y(_03917_)
  );
  OAI21X1 _10352_ (
    .A(_03907_),
    .B(_03909_),
    .C(_03917_),
    .Y(frontend_0.e_state_nxt_0_ )
  );
  AND2X1 _10353_ (
    .A(frontend_0.e_state_nxt_3_ ),
    .B(frontend_0.e_state_nxt_0_ ),
    .Y(_03918_)
  );
  NAND2X1 _10354_ (
    .A(frontend_0.e_state_nxt_3_ ),
    .B(frontend_0.e_state_nxt_0_ ),
    .Y(_03919_)
  );
  AOI21X1 _10355_ (
    .A(_03891_),
    .B(_03896_),
    .C(_03919_),
    .Y(_03920_)
  );
  OAI21X1 _10356_ (
    .A(_03890_),
    .B(_03897_),
    .C(_03918_),
    .Y(_03921_)
  );
  OAI21X1 _10357_ (
    .A(_03863_),
    .B(_03920_),
    .C(_03689_),
    .Y(_03922_)
  );
  NOR3X1 _10358_ (
    .A(_03689_),
    .B(_03863_),
    .C(_03920_),
    .Y(_03923_)
  );
  NAND3X1 _10359_ (
    .A(dbg_0.UNUSED_pc_1_ ),
    .B(_03862_),
    .C(_03921_),
    .Y(_03924_)
  );
  AOI21X1 _10360_ (
    .A(_03922_),
    .B(_03924_),
    .C(frontend_0.i_state_3_ ),
    .Y(_03925_)
  );
  OAI21X1 _10361_ (
    .A(dbg_0.fe_mdb_in_1_ ),
    .B(_03686_),
    .C(_03687_),
    .Y(_03926_)
  );
  OR2X1 _10362_ (
    .A(_03925_),
    .B(_03926_),
    .Y(_03927_)
  );
  OAI21X1 _10363_ (
    .A(execution_unit_0.pc_sw_wr ),
    .B(frontend_0.irq_addr_1_ ),
    .C(_03882_),
    .Y(_03928_)
  );
  AOI21X1 _10364_ (
    .A(_03927_),
    .B(_03928_),
    .C(_03898_),
    .Y(execution_unit_0.pc_nxt_1_ )
  );
  NOR2X1 _10365_ (
    .A(_03683_),
    .B(execution_unit_0.alu_0.alu_out_2_ ),
    .Y(_03929_)
  );
  XNOR2X1 _10366_ (
    .A(_03691_),
    .B(_03923_),
    .Y(_03930_)
  );
  AOI21X1 _10367_ (
    .A(_03678_),
    .B(frontend_0.i_state_3_ ),
    .C(frontend_0.i_state_0_ ),
    .Y(_03931_)
  );
  OAI21X1 _10368_ (
    .A(frontend_0.i_state_3_ ),
    .B(_03930_),
    .C(_03931_),
    .Y(_03932_)
  );
  AOI21X1 _10369_ (
    .A(frontend_0.i_state_0_ ),
    .B(frontend_0.irq_addr_2_ ),
    .C(execution_unit_0.pc_sw_wr ),
    .Y(_03933_)
  );
  AOI21X1 _10370_ (
    .A(_03932_),
    .B(_03933_),
    .C(_03929_),
    .Y(execution_unit_0.pc_nxt_2_ )
  );
  OR2X1 _10371_ (
    .A(_03683_),
    .B(execution_unit_0.alu_0.alu_out_3_ ),
    .Y(_03934_)
  );
  OAI21X1 _10372_ (
    .A(_03691_),
    .B(_03924_),
    .C(_03693_),
    .Y(_03935_)
  );
  NOR3X1 _10373_ (
    .A(_03691_),
    .B(_03693_),
    .C(_03924_),
    .Y(_03936_)
  );
  NAND3X1 _10374_ (
    .A(dbg_0.UNUSED_pc_2_ ),
    .B(dbg_0.UNUSED_pc_3_ ),
    .C(_03923_),
    .Y(_03937_)
  );
  AOI21X1 _10375_ (
    .A(_03935_),
    .B(_03937_),
    .C(frontend_0.i_state_3_ ),
    .Y(_03938_)
  );
  OAI21X1 _10376_ (
    .A(dbg_0.fe_mdb_in_3_ ),
    .B(_03686_),
    .C(_03687_),
    .Y(_03939_)
  );
  OAI21X1 _10377_ (
    .A(execution_unit_0.pc_sw_wr ),
    .B(frontend_0.irq_addr_3_ ),
    .C(_03882_),
    .Y(_03940_)
  );
  OAI21X1 _10378_ (
    .A(_03938_),
    .B(_03939_),
    .C(_03940_),
    .Y(_03941_)
  );
  AND2X1 _10379_ (
    .A(_03934_),
    .B(_03941_),
    .Y(execution_unit_0.pc_nxt_3_ )
  );
  NOR2X1 _10380_ (
    .A(_03683_),
    .B(execution_unit_0.alu_0.alu_out_4_ ),
    .Y(_03942_)
  );
  XNOR2X1 _10381_ (
    .A(_03695_),
    .B(_03936_),
    .Y(_03943_)
  );
  AOI21X1 _10382_ (
    .A(_03675_),
    .B(frontend_0.i_state_3_ ),
    .C(frontend_0.i_state_0_ ),
    .Y(_03944_)
  );
  OAI21X1 _10383_ (
    .A(frontend_0.i_state_3_ ),
    .B(_03943_),
    .C(_03944_),
    .Y(_03945_)
  );
  AOI21X1 _10384_ (
    .A(frontend_0.i_state_0_ ),
    .B(frontend_0.irq_addr_4_ ),
    .C(execution_unit_0.pc_sw_wr ),
    .Y(_03946_)
  );
  AOI21X1 _10385_ (
    .A(_03945_),
    .B(_03946_),
    .C(_03942_),
    .Y(execution_unit_0.pc_nxt_4_ )
  );
  NOR2X1 _10386_ (
    .A(_03683_),
    .B(execution_unit_0.alu_0.alu_out_5_ ),
    .Y(_03947_)
  );
  NOR3X1 _10387_ (
    .A(_03695_),
    .B(_03696_),
    .C(_03937_),
    .Y(_03948_)
  );
  NAND3X1 _10388_ (
    .A(dbg_0.UNUSED_pc_4_ ),
    .B(dbg_0.UNUSED_pc_5_ ),
    .C(_03936_),
    .Y(_03949_)
  );
  OAI21X1 _10389_ (
    .A(_03695_),
    .B(_03937_),
    .C(_03696_),
    .Y(_03950_)
  );
  AOI21X1 _10390_ (
    .A(_03949_),
    .B(_03950_),
    .C(frontend_0.i_state_3_ ),
    .Y(_03951_)
  );
  OAI21X1 _10391_ (
    .A(dbg_0.fe_mdb_in_5_ ),
    .B(_03686_),
    .C(_03687_),
    .Y(_03952_)
  );
  OR2X1 _10392_ (
    .A(_03951_),
    .B(_03952_),
    .Y(_03953_)
  );
  NAND2X1 _10393_ (
    .A(frontend_0.i_state_0_ ),
    .B(frontend_0.irq_addr_5_ ),
    .Y(_03954_)
  );
  AOI21X1 _10394_ (
    .A(frontend_0.i_state_0_ ),
    .B(frontend_0.irq_addr_5_ ),
    .C(execution_unit_0.pc_sw_wr ),
    .Y(_03955_)
  );
  AOI21X1 _10395_ (
    .A(_03953_),
    .B(_03955_),
    .C(_03947_),
    .Y(execution_unit_0.pc_nxt_5_ )
  );
  NOR2X1 _10396_ (
    .A(_03683_),
    .B(execution_unit_0.alu_0.alu_out_6_ ),
    .Y(_03956_)
  );
  XNOR2X1 _10397_ (
    .A(_03697_),
    .B(_03948_),
    .Y(_03957_)
  );
  AOI21X1 _10398_ (
    .A(frontend_0.i_state_3_ ),
    .B(_03698_),
    .C(frontend_0.i_state_0_ ),
    .Y(_03958_)
  );
  OAI21X1 _10399_ (
    .A(frontend_0.i_state_3_ ),
    .B(_03957_),
    .C(_03958_),
    .Y(_03959_)
  );
  AOI21X1 _10400_ (
    .A(frontend_0.i_state_0_ ),
    .B(frontend_0.irq_addr_6_ ),
    .C(execution_unit_0.pc_sw_wr ),
    .Y(_03960_)
  );
  AOI21X1 _10401_ (
    .A(_03959_),
    .B(_03960_),
    .C(_03956_),
    .Y(execution_unit_0.pc_nxt_6_ )
  );
  NOR3X1 _10402_ (
    .A(_03697_),
    .B(_03700_),
    .C(_03949_),
    .Y(_03961_)
  );
  NAND3X1 _10403_ (
    .A(dbg_0.UNUSED_pc_6_ ),
    .B(dbg_0.UNUSED_pc_7_ ),
    .C(_03948_),
    .Y(_03962_)
  );
  OAI21X1 _10404_ (
    .A(_03697_),
    .B(_03949_),
    .C(_03700_),
    .Y(_03963_)
  );
  NAND2X1 _10405_ (
    .A(_03686_),
    .B(_03963_),
    .Y(_03964_)
  );
  AOI21X1 _10406_ (
    .A(dbg_0.fe_mdb_in_7_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03882_),
    .Y(_03965_)
  );
  OAI21X1 _10407_ (
    .A(_03961_),
    .B(_03964_),
    .C(_03965_),
    .Y(_03966_)
  );
  OAI21X1 _10408_ (
    .A(_03683_),
    .B(execution_unit_0.alu_0.alu_out_7_ ),
    .C(_03966_),
    .Y(_03967_)
  );
  INVX1 _10409_ (
    .A(_03967_),
    .Y(execution_unit_0.pc_nxt_7_ )
  );
  NOR2X1 _10410_ (
    .A(_03701_),
    .B(_03962_),
    .Y(_03968_)
  );
  OAI21X1 _10411_ (
    .A(dbg_0.UNUSED_pc_8_ ),
    .B(_03961_),
    .C(_03686_),
    .Y(_03969_)
  );
  AOI21X1 _10412_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03882_),
    .Y(_03970_)
  );
  OAI21X1 _10413_ (
    .A(_03968_),
    .B(_03969_),
    .C(_03970_),
    .Y(_03971_)
  );
  OAI21X1 _10414_ (
    .A(_03683_),
    .B(execution_unit_0.pc_sw_8_ ),
    .C(_03971_),
    .Y(_03972_)
  );
  INVX1 _10415_ (
    .A(_03972_),
    .Y(execution_unit_0.pc_nxt_8_ )
  );
  NOR3X1 _10416_ (
    .A(_03701_),
    .B(_03702_),
    .C(_03962_),
    .Y(_03973_)
  );
  NAND3X1 _10417_ (
    .A(dbg_0.UNUSED_pc_8_ ),
    .B(dbg_0.UNUSED_pc_9_ ),
    .C(_03961_),
    .Y(_03974_)
  );
  OAI21X1 _10418_ (
    .A(_03701_),
    .B(_03962_),
    .C(_03702_),
    .Y(_03975_)
  );
  NAND2X1 _10419_ (
    .A(_03686_),
    .B(_03975_),
    .Y(_03976_)
  );
  AOI21X1 _10420_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03882_),
    .Y(_03977_)
  );
  OAI21X1 _10421_ (
    .A(_03973_),
    .B(_03976_),
    .C(_03977_),
    .Y(_03978_)
  );
  OAI21X1 _10422_ (
    .A(_03683_),
    .B(execution_unit_0.pc_sw_9_ ),
    .C(_03978_),
    .Y(_03979_)
  );
  INVX1 _10423_ (
    .A(_03979_),
    .Y(execution_unit_0.pc_nxt_9_ )
  );
  XNOR2X1 _10424_ (
    .A(dbg_0.UNUSED_pc_10_ ),
    .B(_03973_),
    .Y(_03980_)
  );
  AOI21X1 _10425_ (
    .A(dbg_0.fe_mdb_in_10_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03882_),
    .Y(_03981_)
  );
  OAI21X1 _10426_ (
    .A(frontend_0.i_state_3_ ),
    .B(_03980_),
    .C(_03981_),
    .Y(_03982_)
  );
  OAI21X1 _10427_ (
    .A(_03683_),
    .B(execution_unit_0.pc_sw_10_ ),
    .C(_03982_),
    .Y(_03983_)
  );
  INVX1 _10428_ (
    .A(_03983_),
    .Y(execution_unit_0.pc_nxt_10_ )
  );
  NOR3X1 _10429_ (
    .A(_03703_),
    .B(_03704_),
    .C(_03974_),
    .Y(_03984_)
  );
  NAND3X1 _10430_ (
    .A(dbg_0.UNUSED_pc_10_ ),
    .B(dbg_0.UNUSED_pc_11_ ),
    .C(_03973_),
    .Y(_03985_)
  );
  OAI21X1 _10431_ (
    .A(_03703_),
    .B(_03974_),
    .C(_03704_),
    .Y(_03986_)
  );
  NAND2X1 _10432_ (
    .A(_03686_),
    .B(_03986_),
    .Y(_03987_)
  );
  AOI21X1 _10433_ (
    .A(dbg_0.fe_mdb_in_11_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03882_),
    .Y(_03988_)
  );
  OAI21X1 _10434_ (
    .A(_03984_),
    .B(_03987_),
    .C(_03988_),
    .Y(_03989_)
  );
  OAI21X1 _10435_ (
    .A(_03683_),
    .B(execution_unit_0.pc_sw_11_ ),
    .C(_03989_),
    .Y(_03990_)
  );
  INVX1 _10436_ (
    .A(_03990_),
    .Y(execution_unit_0.pc_nxt_11_ )
  );
  NOR2X1 _10437_ (
    .A(_03683_),
    .B(execution_unit_0.pc_sw_12_ ),
    .Y(_03991_)
  );
  AOI21X1 _10438_ (
    .A(_03705_),
    .B(_03985_),
    .C(frontend_0.i_state_3_ ),
    .Y(_03992_)
  );
  OAI21X1 _10439_ (
    .A(_03705_),
    .B(_03985_),
    .C(_03992_),
    .Y(_03993_)
  );
  AOI21X1 _10440_ (
    .A(frontend_0.i_state_3_ ),
    .B(dbg_0.fe_mdb_in_12_ ),
    .C(_03882_),
    .Y(_03994_)
  );
  AOI21X1 _10441_ (
    .A(_03993_),
    .B(_03994_),
    .C(_03991_),
    .Y(execution_unit_0.pc_nxt_12_ )
  );
  NOR2X1 _10442_ (
    .A(_03683_),
    .B(execution_unit_0.pc_sw_13_ ),
    .Y(_03995_)
  );
  NOR3X1 _10443_ (
    .A(_03705_),
    .B(_03707_),
    .C(_03985_),
    .Y(_03996_)
  );
  NAND3X1 _10444_ (
    .A(dbg_0.UNUSED_pc_12_ ),
    .B(dbg_0.UNUSED_pc_13_ ),
    .C(_03984_),
    .Y(_03997_)
  );
  OAI21X1 _10445_ (
    .A(_03705_),
    .B(_03985_),
    .C(_03707_),
    .Y(_03998_)
  );
  NAND3X1 _10446_ (
    .A(_03686_),
    .B(_03997_),
    .C(_03998_),
    .Y(_03999_)
  );
  AOI21X1 _10447_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03882_),
    .Y(_04000_)
  );
  AOI21X1 _10448_ (
    .A(_03999_),
    .B(_04000_),
    .C(_03995_),
    .Y(execution_unit_0.pc_nxt_13_ )
  );
  NOR2X1 _10449_ (
    .A(_03683_),
    .B(execution_unit_0.pc_sw_14_ ),
    .Y(_04001_)
  );
  AOI21X1 _10450_ (
    .A(_03708_),
    .B(_03997_),
    .C(frontend_0.i_state_3_ ),
    .Y(_04002_)
  );
  OAI21X1 _10451_ (
    .A(_03708_),
    .B(_03997_),
    .C(_04002_),
    .Y(_04003_)
  );
  AOI21X1 _10452_ (
    .A(dbg_0.fe_mdb_in_14_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03882_),
    .Y(_04004_)
  );
  AOI21X1 _10453_ (
    .A(_04003_),
    .B(_04004_),
    .C(_04001_),
    .Y(execution_unit_0.pc_nxt_14_ )
  );
  NOR2X1 _10454_ (
    .A(_03683_),
    .B(execution_unit_0.pc_sw_15_ ),
    .Y(_04005_)
  );
  OAI21X1 _10455_ (
    .A(_03708_),
    .B(_03997_),
    .C(_03709_),
    .Y(_04006_)
  );
  NAND3X1 _10456_ (
    .A(dbg_0.UNUSED_pc_14_ ),
    .B(dbg_0.UNUSED_pc_15_ ),
    .C(_03996_),
    .Y(_04007_)
  );
  NAND3X1 _10457_ (
    .A(_03686_),
    .B(_04006_),
    .C(_04007_),
    .Y(_04008_)
  );
  AOI21X1 _10458_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03882_),
    .Y(_04009_)
  );
  AOI21X1 _10459_ (
    .A(_04008_),
    .B(_04009_),
    .C(_04005_),
    .Y(execution_unit_0.pc_nxt_15_ )
  );
  NOR2X1 _10460_ (
    .A(frontend_0.inst_dest_bin_3_ ),
    .B(frontend_0.inst_dest_bin_2_ ),
    .Y(_04010_)
  );
  NOR2X1 _10461_ (
    .A(frontend_0.inst_dest_bin_0_ ),
    .B(frontend_0.inst_dest_bin_1_ ),
    .Y(_04011_)
  );
  AND2X1 _10462_ (
    .A(_04010_),
    .B(_04011_),
    .Y(_04012_)
  );
  NOR2X1 _10463_ (
    .A(execution_unit_0.alu_0.inst_so_7_ ),
    .B(_03840_),
    .Y(_04013_)
  );
  INVX1 _10464_ (
    .A(_04013_),
    .Y(_04014_)
  );
  AOI21X1 _10465_ (
    .A(_04012_),
    .B(_04013_),
    .C(execution_unit_0.inst_type_1_ ),
    .Y(_04015_)
  );
  NAND2X1 _10466_ (
    .A(_03715_),
    .B(_03716_),
    .Y(_04016_)
  );
  NAND3X1 _10467_ (
    .A(cpu_halt_st),
    .B(_03717_),
    .C(_03718_),
    .Y(_04017_)
  );
  OAI22X1 _10468_ (
    .A(cpu_halt_st),
    .B(_04015_),
    .C(_04016_),
    .D(_04017_),
    .Y(execution_unit_0.inst_dest_0_ )
  );
  NOR2X1 _10469_ (
    .A(_03712_),
    .B(frontend_0.inst_dest_bin_1_ ),
    .Y(_04018_)
  );
  AND2X1 _10470_ (
    .A(_04010_),
    .B(_04018_),
    .Y(_04019_)
  );
  NOR2X1 _10471_ (
    .A(cpu_halt_st),
    .B(execution_unit_0.inst_type_1_ ),
    .Y(_04020_)
  );
  OAI21X1 _10472_ (
    .A(_04014_),
    .B(_04019_),
    .C(_04020_),
    .Y(_04021_)
  );
  NAND2X1 _10473_ (
    .A(dbg_0.dbg_mem_addr_0_ ),
    .B(_03716_),
    .Y(_04022_)
  );
  OAI21X1 _10474_ (
    .A(_04017_),
    .B(_04022_),
    .C(_04021_),
    .Y(execution_unit_0.inst_dest_1_ )
  );
  NOR2X1 _10475_ (
    .A(frontend_0.inst_dest_bin_0_ ),
    .B(_03713_),
    .Y(_04023_)
  );
  NAND2X1 _10476_ (
    .A(_04010_),
    .B(_04023_),
    .Y(_04024_)
  );
  NAND2X1 _10477_ (
    .A(_04013_),
    .B(_04020_),
    .Y(_04025_)
  );
  NAND2X1 _10478_ (
    .A(_03715_),
    .B(dbg_0.dbg_mem_addr_1_ ),
    .Y(_04026_)
  );
  OAI22X1 _10479_ (
    .A(_04024_),
    .B(_04025_),
    .C(_04026_),
    .D(_04017_),
    .Y(execution_unit_0.inst_dest_2_ )
  );
  NOR2X1 _10480_ (
    .A(_03712_),
    .B(_03713_),
    .Y(_04027_)
  );
  NAND2X1 _10481_ (
    .A(_04010_),
    .B(_04027_),
    .Y(_04028_)
  );
  NAND2X1 _10482_ (
    .A(dbg_0.dbg_mem_addr_0_ ),
    .B(dbg_0.dbg_mem_addr_1_ ),
    .Y(_04029_)
  );
  OAI22X1 _10483_ (
    .A(_04025_),
    .B(_04028_),
    .C(_04029_),
    .D(_04017_),
    .Y(execution_unit_0.inst_dest_3_ )
  );
  NOR2X1 _10484_ (
    .A(frontend_0.inst_dest_bin_3_ ),
    .B(_03711_),
    .Y(_04030_)
  );
  NAND2X1 _10485_ (
    .A(_04011_),
    .B(_04030_),
    .Y(_04031_)
  );
  NAND2X1 _10486_ (
    .A(_03717_),
    .B(dbg_0.dbg_mem_addr_2_ ),
    .Y(_04032_)
  );
  NAND3X1 _10487_ (
    .A(cpu_halt_st),
    .B(_03715_),
    .C(_03716_),
    .Y(_04033_)
  );
  OAI22X1 _10488_ (
    .A(_04025_),
    .B(_04031_),
    .C(_04032_),
    .D(_04033_),
    .Y(execution_unit_0.inst_dest_4_ )
  );
  NAND2X1 _10489_ (
    .A(_04018_),
    .B(_04030_),
    .Y(_04034_)
  );
  NAND3X1 _10490_ (
    .A(cpu_halt_st),
    .B(dbg_0.dbg_mem_addr_0_ ),
    .C(_03716_),
    .Y(_04035_)
  );
  OAI22X1 _10491_ (
    .A(_04025_),
    .B(_04034_),
    .C(_04035_),
    .D(_04032_),
    .Y(execution_unit_0.inst_dest_5_ )
  );
  NAND2X1 _10492_ (
    .A(_04023_),
    .B(_04030_),
    .Y(_04036_)
  );
  NAND3X1 _10493_ (
    .A(cpu_halt_st),
    .B(_03715_),
    .C(dbg_0.dbg_mem_addr_1_ ),
    .Y(_04037_)
  );
  OAI22X1 _10494_ (
    .A(_04025_),
    .B(_04036_),
    .C(_04037_),
    .D(_04032_),
    .Y(execution_unit_0.inst_dest_6_ )
  );
  NAND2X1 _10495_ (
    .A(_04027_),
    .B(_04030_),
    .Y(_04038_)
  );
  NAND3X1 _10496_ (
    .A(cpu_halt_st),
    .B(dbg_0.dbg_mem_addr_0_ ),
    .C(dbg_0.dbg_mem_addr_1_ ),
    .Y(_04039_)
  );
  OAI22X1 _10497_ (
    .A(_04025_),
    .B(_04038_),
    .C(_04039_),
    .D(_04032_),
    .Y(execution_unit_0.inst_dest_7_ )
  );
  NOR2X1 _10498_ (
    .A(_03710_),
    .B(frontend_0.inst_dest_bin_2_ ),
    .Y(_04040_)
  );
  NAND2X1 _10499_ (
    .A(_04011_),
    .B(_04040_),
    .Y(_04041_)
  );
  NAND2X1 _10500_ (
    .A(dbg_0.dbg_mem_addr_3_ ),
    .B(_03718_),
    .Y(_04042_)
  );
  OAI22X1 _10501_ (
    .A(_04025_),
    .B(_04041_),
    .C(_04042_),
    .D(_04033_),
    .Y(execution_unit_0.inst_dest_8_ )
  );
  NAND2X1 _10502_ (
    .A(_04018_),
    .B(_04040_),
    .Y(_04043_)
  );
  OAI22X1 _10503_ (
    .A(_04035_),
    .B(_04042_),
    .C(_04043_),
    .D(_04025_),
    .Y(execution_unit_0.inst_dest_9_ )
  );
  NAND2X1 _10504_ (
    .A(_04023_),
    .B(_04040_),
    .Y(_04044_)
  );
  OAI22X1 _10505_ (
    .A(_04037_),
    .B(_04042_),
    .C(_04044_),
    .D(_04025_),
    .Y(execution_unit_0.inst_dest_10_ )
  );
  NAND2X1 _10506_ (
    .A(_04027_),
    .B(_04040_),
    .Y(_04045_)
  );
  OAI22X1 _10507_ (
    .A(_04039_),
    .B(_04042_),
    .C(_04045_),
    .D(_04025_),
    .Y(execution_unit_0.inst_dest_11_ )
  );
  NOR2X1 _10508_ (
    .A(_03710_),
    .B(_03711_),
    .Y(_04046_)
  );
  NAND2X1 _10509_ (
    .A(_04011_),
    .B(_04046_),
    .Y(_04047_)
  );
  NAND2X1 _10510_ (
    .A(dbg_0.dbg_mem_addr_3_ ),
    .B(dbg_0.dbg_mem_addr_2_ ),
    .Y(_04048_)
  );
  OAI22X1 _10511_ (
    .A(_04025_),
    .B(_04047_),
    .C(_04048_),
    .D(_04033_),
    .Y(execution_unit_0.inst_dest_12_ )
  );
  NAND2X1 _10512_ (
    .A(_04018_),
    .B(_04046_),
    .Y(_04049_)
  );
  OAI22X1 _10513_ (
    .A(_04035_),
    .B(_04048_),
    .C(_04049_),
    .D(_04025_),
    .Y(execution_unit_0.inst_dest_13_ )
  );
  NAND2X1 _10514_ (
    .A(_04023_),
    .B(_04046_),
    .Y(_04050_)
  );
  OAI22X1 _10515_ (
    .A(_04037_),
    .B(_04048_),
    .C(_04050_),
    .D(_04025_),
    .Y(execution_unit_0.inst_dest_14_ )
  );
  NAND2X1 _10516_ (
    .A(_04027_),
    .B(_04046_),
    .Y(_04051_)
  );
  OAI22X1 _10517_ (
    .A(_04039_),
    .B(_04048_),
    .C(_04051_),
    .D(_04025_),
    .Y(execution_unit_0.inst_dest_15_ )
  );
  AND2X1 _10518_ (
    .A(execution_unit_0.inst_type_0_ ),
    .B(_04012_),
    .Y(_04052_)
  );
  NOR2X1 _10519_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(execution_unit_0.inst_type_2_ ),
    .Y(_04053_)
  );
  OAI21X1 _10520_ (
    .A(execution_unit_0.alu_0.inst_so_7_ ),
    .B(_04052_),
    .C(_04053_),
    .Y(_04054_)
  );
  OR2X1 _10521_ (
    .A(frontend_0.inst_src_bin_0_ ),
    .B(frontend_0.inst_src_bin_1_ ),
    .Y(_04055_)
  );
  NAND3X1 _10522_ (
    .A(_03721_),
    .B(_03722_),
    .C(execution_unit_0.inst_type_2_ ),
    .Y(_04056_)
  );
  OAI21X1 _10523_ (
    .A(_04055_),
    .B(_04056_),
    .C(_04054_),
    .Y(execution_unit_0.inst_src_0_ )
  );
  NOR2X1 _10524_ (
    .A(execution_unit_0.alu_0.inst_so_7_ ),
    .B(_03719_),
    .Y(_04057_)
  );
  AOI21X1 _10525_ (
    .A(_04019_),
    .B(_04057_),
    .C(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .Y(_04058_)
  );
  NAND2X1 _10526_ (
    .A(frontend_0.inst_src_bin_0_ ),
    .B(_03720_),
    .Y(_04059_)
  );
  OAI22X1 _10527_ (
    .A(execution_unit_0.inst_type_2_ ),
    .B(_04058_),
    .C(_04059_),
    .D(_04056_),
    .Y(execution_unit_0.inst_src_1_ )
  );
  NAND2X1 _10528_ (
    .A(_04053_),
    .B(_04057_),
    .Y(_04060_)
  );
  OR2X1 _10529_ (
    .A(frontend_0.inst_src_bin_0_ ),
    .B(_03720_),
    .Y(_04061_)
  );
  OAI22X1 _10530_ (
    .A(_04024_),
    .B(_04060_),
    .C(_04061_),
    .D(_04056_),
    .Y(execution_unit_0.inst_src_2_ )
  );
  NAND2X1 _10531_ (
    .A(frontend_0.inst_src_bin_0_ ),
    .B(frontend_0.inst_src_bin_1_ ),
    .Y(_04062_)
  );
  OAI22X1 _10532_ (
    .A(_04028_),
    .B(_04060_),
    .C(_04062_),
    .D(_04056_),
    .Y(execution_unit_0.inst_src_3_ )
  );
  NAND2X1 _10533_ (
    .A(_03721_),
    .B(frontend_0.inst_src_bin_2_ ),
    .Y(_04063_)
  );
  OR2X1 _10534_ (
    .A(_03723_),
    .B(_04055_),
    .Y(_04064_)
  );
  OAI22X1 _10535_ (
    .A(_04031_),
    .B(_04060_),
    .C(_04063_),
    .D(_04064_),
    .Y(execution_unit_0.inst_src_4_ )
  );
  OR2X1 _10536_ (
    .A(_03723_),
    .B(_04059_),
    .Y(_04065_)
  );
  OAI22X1 _10537_ (
    .A(_04034_),
    .B(_04060_),
    .C(_04063_),
    .D(_04065_),
    .Y(execution_unit_0.inst_src_5_ )
  );
  OR2X1 _10538_ (
    .A(_03723_),
    .B(_04061_),
    .Y(_04066_)
  );
  OAI22X1 _10539_ (
    .A(_04036_),
    .B(_04060_),
    .C(_04063_),
    .D(_04066_),
    .Y(execution_unit_0.inst_src_6_ )
  );
  OR2X1 _10540_ (
    .A(_03723_),
    .B(_04062_),
    .Y(_04067_)
  );
  OAI22X1 _10541_ (
    .A(_04038_),
    .B(_04060_),
    .C(_04063_),
    .D(_04067_),
    .Y(execution_unit_0.inst_src_7_ )
  );
  NAND2X1 _10542_ (
    .A(frontend_0.inst_src_bin_3_ ),
    .B(_03722_),
    .Y(_04068_)
  );
  OAI22X1 _10543_ (
    .A(_04041_),
    .B(_04060_),
    .C(_04064_),
    .D(_04068_),
    .Y(execution_unit_0.inst_src_8_ )
  );
  OAI22X1 _10544_ (
    .A(_04043_),
    .B(_04060_),
    .C(_04065_),
    .D(_04068_),
    .Y(execution_unit_0.inst_src_9_ )
  );
  OAI22X1 _10545_ (
    .A(_04044_),
    .B(_04060_),
    .C(_04066_),
    .D(_04068_),
    .Y(execution_unit_0.inst_src_10_ )
  );
  OAI22X1 _10546_ (
    .A(_04045_),
    .B(_04060_),
    .C(_04067_),
    .D(_04068_),
    .Y(execution_unit_0.inst_src_11_ )
  );
  NAND2X1 _10547_ (
    .A(frontend_0.inst_src_bin_3_ ),
    .B(frontend_0.inst_src_bin_2_ ),
    .Y(_04069_)
  );
  OAI22X1 _10548_ (
    .A(_04047_),
    .B(_04060_),
    .C(_04064_),
    .D(_04069_),
    .Y(execution_unit_0.inst_src_12_ )
  );
  OAI22X1 _10549_ (
    .A(_04049_),
    .B(_04060_),
    .C(_04065_),
    .D(_04069_),
    .Y(execution_unit_0.inst_src_13_ )
  );
  OAI22X1 _10550_ (
    .A(_04050_),
    .B(_04060_),
    .C(_04066_),
    .D(_04069_),
    .Y(execution_unit_0.inst_src_14_ )
  );
  OAI22X1 _10551_ (
    .A(_04051_),
    .B(_04060_),
    .C(_04067_),
    .D(_04069_),
    .Y(execution_unit_0.inst_src_15_ )
  );
  NOR2X1 _10552_ (
    .A(_03766_),
    .B(dbg_0.decode_noirq ),
    .Y(_04070_)
  );
  OAI21X1 _10553_ (
    .A(_03682_),
    .B(_03861_),
    .C(_03767_),
    .Y(_04071_)
  );
  AND2X1 _10554_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(_03767_),
    .Y(_04072_)
  );
  OAI21X1 _10555_ (
    .A(_03749_),
    .B(_03765_),
    .C(dbg_0.fe_mdb_in_15_ ),
    .Y(_04073_)
  );
  NAND2X1 _10556_ (
    .A(_03674_),
    .B(_04072_),
    .Y(_04074_)
  );
  NOR2X1 _10557_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(dbg_0.fe_mdb_in_12_ ),
    .Y(_04075_)
  );
  OAI21X1 _10558_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(_04074_),
    .C(_04071_),
    .Y(_04076_)
  );
  NAND2X1 _10559_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(dbg_0.fe_mdb_in_12_ ),
    .Y(_04077_)
  );
  NOR2X1 _10560_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(_03674_),
    .Y(_04078_)
  );
  AND2X1 _10561_ (
    .A(_03767_),
    .B(_04078_),
    .Y(_04079_)
  );
  INVX1 _10562_ (
    .A(_04079_),
    .Y(_04080_)
  );
  NAND2X1 _10563_ (
    .A(dbg_0.fe_mdb_in_14_ ),
    .B(_04072_),
    .Y(_04081_)
  );
  NAND3X1 _10564_ (
    .A(dbg_0.fe_mdb_in_14_ ),
    .B(_04072_),
    .C(_04075_),
    .Y(_04082_)
  );
  OAI21X1 _10565_ (
    .A(_04077_),
    .B(_04080_),
    .C(_04082_),
    .Y(_04083_)
  );
  OAI22X1 _10566_ (
    .A(execution_unit_0.alu_0.inst_alu_0_ ),
    .B(_04071_),
    .C(_04076_),
    .D(_04083_),
    .Y(_04084_)
  );
  INVX1 _10567_ (
    .A(_04084_),
    .Y(_03349_)
  );
  OAI21X1 _10568_ (
    .A(execution_unit_0.alu_0.inst_alu_1_ ),
    .B(_04071_),
    .C(_04076_),
    .Y(_04085_)
  );
  INVX1 _10569_ (
    .A(_04085_),
    .Y(_03351_)
  );
  NAND2X1 _10570_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(dbg_0.decode_noirq ),
    .Y(_04086_)
  );
  OR2X1 _10571_ (
    .A(dbg_0.fe_mdb_in_12_ ),
    .B(_04086_),
    .Y(_04087_)
  );
  OR2X1 _10572_ (
    .A(_04074_),
    .B(_04087_),
    .Y(_04088_)
  );
  OAI21X1 _10573_ (
    .A(_04080_),
    .B(_04086_),
    .C(_04088_),
    .Y(_04089_)
  );
  AOI21X1 _10574_ (
    .A(execution_unit_0.alu_0.inst_alu_2_ ),
    .B(_04070_),
    .C(_04089_),
    .Y(_04090_)
  );
  INVX1 _10575_ (
    .A(_04090_),
    .Y(_03352_)
  );
  OAI21X1 _10576_ (
    .A(_03673_),
    .B(_03769_),
    .C(_03798_),
    .Y(_04091_)
  );
  OAI22X1 _10577_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(_04074_),
    .C(_04075_),
    .D(_04080_),
    .Y(_04092_)
  );
  OAI21X1 _10578_ (
    .A(_04091_),
    .B(_04092_),
    .C(_04071_),
    .Y(_04093_)
  );
  OAI21X1 _10579_ (
    .A(_03724_),
    .B(_04071_),
    .C(_04093_),
    .Y(_03353_)
  );
  NOR2X1 _10580_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_04071_),
    .Y(_04094_)
  );
  NOR2X1 _10581_ (
    .A(_04073_),
    .B(_04077_),
    .Y(_04095_)
  );
  NOR2X1 _10582_ (
    .A(_04070_),
    .B(_04095_),
    .Y(_04096_)
  );
  AOI21X1 _10583_ (
    .A(_04082_),
    .B(_04096_),
    .C(_04094_),
    .Y(_03354_)
  );
  NAND2X1 _10584_ (
    .A(execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_04070_),
    .Y(_04097_)
  );
  NAND2X1 _10585_ (
    .A(_03806_),
    .B(dbg_0.decode_noirq ),
    .Y(_04098_)
  );
  NOR2X1 _10586_ (
    .A(_03674_),
    .B(_03706_),
    .Y(_04099_)
  );
  NAND3X1 _10587_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(_03673_),
    .C(_04099_),
    .Y(_04100_)
  );
  OAI21X1 _10588_ (
    .A(_04098_),
    .B(_04100_),
    .C(_04097_),
    .Y(_03355_)
  );
  NAND2X1 _10589_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_04070_),
    .Y(_04101_)
  );
  OAI21X1 _10590_ (
    .A(_04081_),
    .B(_04087_),
    .C(_04101_),
    .Y(_03356_)
  );
  OAI21X1 _10591_ (
    .A(_03725_),
    .B(_04071_),
    .C(_04088_),
    .Y(_03357_)
  );
  NOR2X1 _10592_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(_03774_),
    .Y(_04102_)
  );
  OAI21X1 _10593_ (
    .A(_04095_),
    .B(_04102_),
    .C(_04071_),
    .Y(_04103_)
  );
  OAI21X1 _10594_ (
    .A(_03726_),
    .B(_04071_),
    .C(_04103_),
    .Y(_03358_)
  );
  NOR2X1 _10595_ (
    .A(execution_unit_0.alu_0.inst_alu_9_ ),
    .B(_04071_),
    .Y(_04104_)
  );
  AOI21X1 _10596_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(_04072_),
    .C(_04092_),
    .Y(_04105_)
  );
  NOR2X1 _10597_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(dbg_0.fe_mdb_in_7_ ),
    .Y(_04106_)
  );
  INVX1 _10598_ (
    .A(_04106_),
    .Y(_04107_)
  );
  AOI21X1 _10599_ (
    .A(_03770_),
    .B(_04106_),
    .C(_04070_),
    .Y(_04108_)
  );
  OAI21X1 _10600_ (
    .A(_03771_),
    .B(_04107_),
    .C(_04071_),
    .Y(_04109_)
  );
  NOR2X1 _10601_ (
    .A(_04102_),
    .B(_04109_),
    .Y(_04110_)
  );
  AOI21X1 _10602_ (
    .A(_04105_),
    .B(_04110_),
    .C(_04104_),
    .Y(_03359_)
  );
  OAI21X1 _10603_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(_04071_),
    .C(_04109_),
    .Y(_04111_)
  );
  INVX1 _10604_ (
    .A(_04111_),
    .Y(_03350_)
  );
  NAND2X1 _10605_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_alu ),
    .B(_04070_),
    .Y(_04112_)
  );
  NAND3X1 _10606_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(_03674_),
    .C(dbg_0.fe_mdb_in_12_ ),
    .Y(_04113_)
  );
  OAI21X1 _10607_ (
    .A(_04098_),
    .B(_04113_),
    .C(_04112_),
    .Y(_03437_)
  );
  NOR2X1 _10608_ (
    .A(_03829_),
    .B(_03912_),
    .Y(_03341_)
  );
  NAND2X1 _10609_ (
    .A(execution_unit_0.inst_ad_0_ ),
    .B(_04070_),
    .Y(_04114_)
  );
  OAI21X1 _10610_ (
    .A(dbg_0.fe_mdb_in_7_ ),
    .B(_04098_),
    .C(_04114_),
    .Y(_03345_)
  );
  OR2X1 _10611_ (
    .A(_03672_),
    .B(_04098_),
    .Y(_04115_)
  );
  NOR2X1 _10612_ (
    .A(dbg_0.fe_mdb_in_0_ ),
    .B(_03784_),
    .Y(_04116_)
  );
  OAI22X1 _10613_ (
    .A(_03680_),
    .B(_04071_),
    .C(_04115_),
    .D(_04116_),
    .Y(_03346_)
  );
  NAND2X1 _10614_ (
    .A(execution_unit_0.UNUSED_inst_ad_symb ),
    .B(_04070_),
    .Y(_04117_)
  );
  NAND2X1 _10615_ (
    .A(_03677_),
    .B(_04116_),
    .Y(_04118_)
  );
  OAI21X1 _10616_ (
    .A(_04115_),
    .B(_04118_),
    .C(_04117_),
    .Y(_03347_)
  );
  NAND2X1 _10617_ (
    .A(execution_unit_0.inst_ad_6_ ),
    .B(_04070_),
    .Y(_04119_)
  );
  NAND2X1 _10618_ (
    .A(dbg_0.fe_mdb_in_1_ ),
    .B(_04116_),
    .Y(_04120_)
  );
  OAI21X1 _10619_ (
    .A(_04115_),
    .B(_04120_),
    .C(_04119_),
    .Y(_03348_)
  );
  OAI21X1 _10620_ (
    .A(_03807_),
    .B(_03875_),
    .C(_04071_),
    .Y(_04121_)
  );
  OAI22X1 _10621_ (
    .A(_03684_),
    .B(_04071_),
    .C(_04121_),
    .D(_03876_),
    .Y(_03421_)
  );
  OAI21X1 _10622_ (
    .A(frontend_0.inst_sz_1_ ),
    .B(_04071_),
    .C(_04121_),
    .Y(_04122_)
  );
  INVX1 _10623_ (
    .A(_04122_),
    .Y(_03422_)
  );
  NAND2X1 _10624_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(_04070_),
    .Y(_04123_)
  );
  NOR2X1 _10625_ (
    .A(_03698_),
    .B(_03766_),
    .Y(_04124_)
  );
  NAND3X1 _10626_ (
    .A(_03778_),
    .B(dbg_0.decode_noirq ),
    .C(_04124_),
    .Y(_04125_)
  );
  OAI21X1 _10627_ (
    .A(_03762_),
    .B(_04125_),
    .C(_04123_),
    .Y(_03368_)
  );
  NOR2X1 _10628_ (
    .A(dbg_0.fe_mdb_in_4_ ),
    .B(dbg_0.fe_mdb_in_5_ ),
    .Y(_04126_)
  );
  NOR2X1 _10629_ (
    .A(execution_unit_0.inst_as_0_ ),
    .B(_04071_),
    .Y(_04127_)
  );
  AOI21X1 _10630_ (
    .A(_03815_),
    .B(_04126_),
    .C(_04070_),
    .Y(_04128_)
  );
  AOI21X1 _10631_ (
    .A(_03778_),
    .B(_04128_),
    .C(_04127_),
    .Y(_03360_)
  );
  OAI21X1 _10632_ (
    .A(_03766_),
    .B(dbg_0.decode_noirq ),
    .C(_03817_),
    .Y(_04129_)
  );
  NOR2X1 _10633_ (
    .A(_03791_),
    .B(_04129_),
    .Y(_04130_)
  );
  AOI22X1 _10634_ (
    .A(execution_unit_0.inst_as_1_ ),
    .B(_04070_),
    .C(_04130_),
    .D(_03801_),
    .Y(_04131_)
  );
  INVX1 _10635_ (
    .A(_04131_),
    .Y(_03361_)
  );
  OAI21X1 _10636_ (
    .A(_03791_),
    .B(_03794_),
    .C(_04071_),
    .Y(_04132_)
  );
  OAI21X1 _10637_ (
    .A(execution_unit_0.inst_as_2_ ),
    .B(_04071_),
    .C(_04132_),
    .Y(_04133_)
  );
  INVX1 _10638_ (
    .A(_04133_),
    .Y(_03362_)
  );
  NAND2X1 _10639_ (
    .A(execution_unit_0.inst_as_3_ ),
    .B(_04070_),
    .Y(_04134_)
  );
  OAI21X1 _10640_ (
    .A(_03802_),
    .B(_04070_),
    .C(_04134_),
    .Y(_03363_)
  );
  NAND2X1 _10641_ (
    .A(execution_unit_0.inst_as_4_ ),
    .B(_04070_),
    .Y(_04135_)
  );
  OAI21X1 _10642_ (
    .A(_03801_),
    .B(_04129_),
    .C(_04135_),
    .Y(_03364_)
  );
  NAND2X1 _10643_ (
    .A(execution_unit_0.inst_as_5_ ),
    .B(_04070_),
    .Y(_04136_)
  );
  OAI21X1 _10644_ (
    .A(_03803_),
    .B(_04070_),
    .C(_04136_),
    .Y(_03365_)
  );
  NAND2X1 _10645_ (
    .A(_03791_),
    .B(_03800_),
    .Y(_04137_)
  );
  NAND2X1 _10646_ (
    .A(execution_unit_0.inst_as_6_ ),
    .B(_04070_),
    .Y(_04138_)
  );
  OAI21X1 _10647_ (
    .A(_04129_),
    .B(_04137_),
    .C(_04138_),
    .Y(_03366_)
  );
  OAI21X1 _10648_ (
    .A(_03673_),
    .B(_03769_),
    .C(_03814_),
    .Y(_04139_)
  );
  OAI21X1 _10649_ (
    .A(_03781_),
    .B(_04137_),
    .C(_04139_),
    .Y(_04140_)
  );
  AND2X1 _10650_ (
    .A(_04071_),
    .B(_04140_),
    .Y(_04141_)
  );
  AOI21X1 _10651_ (
    .A(execution_unit_0.inst_as_7_ ),
    .B(_04070_),
    .C(_04141_),
    .Y(_04142_)
  );
  INVX1 _10652_ (
    .A(_04142_),
    .Y(_03367_)
  );
  NAND2X1 _10653_ (
    .A(execution_unit_0.inst_mov ),
    .B(_04070_),
    .Y(_04143_)
  );
  NAND2X1 _10654_ (
    .A(_04075_),
    .B(_04078_),
    .Y(_04144_)
  );
  OAI21X1 _10655_ (
    .A(_04098_),
    .B(_04144_),
    .C(_04143_),
    .Y(_03393_)
  );
  OAI21X1 _10656_ (
    .A(_03766_),
    .B(dbg_0.decode_noirq ),
    .C(_03671_),
    .Y(_04145_)
  );
  OAI21X1 _10657_ (
    .A(frontend_0.inst_src_bin_0_ ),
    .B(_04071_),
    .C(_04145_),
    .Y(_04146_)
  );
  INVX1 _10658_ (
    .A(_04146_),
    .Y(_03417_)
  );
  OAI21X1 _10659_ (
    .A(_03766_),
    .B(dbg_0.decode_noirq ),
    .C(_03670_),
    .Y(_04147_)
  );
  OAI21X1 _10660_ (
    .A(frontend_0.inst_src_bin_1_ ),
    .B(_04071_),
    .C(_04147_),
    .Y(_04148_)
  );
  INVX1 _10661_ (
    .A(_04148_),
    .Y(_03418_)
  );
  OAI21X1 _10662_ (
    .A(_03766_),
    .B(dbg_0.decode_noirq ),
    .C(dbg_0.fe_mdb_in_10_ ),
    .Y(_04149_)
  );
  OAI21X1 _10663_ (
    .A(_03722_),
    .B(_04071_),
    .C(_04149_),
    .Y(_03419_)
  );
  OAI21X1 _10664_ (
    .A(_03766_),
    .B(dbg_0.decode_noirq ),
    .C(dbg_0.fe_mdb_in_11_ ),
    .Y(_04150_)
  );
  OAI21X1 _10665_ (
    .A(_03721_),
    .B(_04071_),
    .C(_04150_),
    .Y(_03420_)
  );
  OAI21X1 _10666_ (
    .A(_03766_),
    .B(dbg_0.decode_noirq ),
    .C(dbg_0.fe_mdb_in_0_ ),
    .Y(_04151_)
  );
  OAI21X1 _10667_ (
    .A(_03712_),
    .B(_04071_),
    .C(_04151_),
    .Y(_03369_)
  );
  OAI21X1 _10668_ (
    .A(_03766_),
    .B(dbg_0.decode_noirq ),
    .C(dbg_0.fe_mdb_in_1_ ),
    .Y(_04152_)
  );
  OAI21X1 _10669_ (
    .A(_03713_),
    .B(_04071_),
    .C(_04152_),
    .Y(_03370_)
  );
  OAI21X1 _10670_ (
    .A(_03766_),
    .B(dbg_0.decode_noirq ),
    .C(dbg_0.fe_mdb_in_2_ ),
    .Y(_04153_)
  );
  OAI21X1 _10671_ (
    .A(_03711_),
    .B(_04071_),
    .C(_04153_),
    .Y(_03371_)
  );
  OAI21X1 _10672_ (
    .A(_03766_),
    .B(dbg_0.decode_noirq ),
    .C(dbg_0.fe_mdb_in_3_ ),
    .Y(_04154_)
  );
  OAI21X1 _10673_ (
    .A(_03710_),
    .B(_04071_),
    .C(_04154_),
    .Y(_03372_)
  );
  NAND2X1 _10674_ (
    .A(_03770_),
    .B(dbg_0.decode_noirq ),
    .Y(_04155_)
  );
  OAI21X1 _10675_ (
    .A(_03719_),
    .B(_04071_),
    .C(_04155_),
    .Y(_03423_)
  );
  AND2X1 _10676_ (
    .A(_03779_),
    .B(dbg_0.decode_noirq ),
    .Y(_04156_)
  );
  NAND2X1 _10677_ (
    .A(_03779_),
    .B(dbg_0.decode_noirq ),
    .Y(_04157_)
  );
  OAI21X1 _10678_ (
    .A(_03714_),
    .B(_04071_),
    .C(_04157_),
    .Y(_03424_)
  );
  OAI21X1 _10679_ (
    .A(_03723_),
    .B(_04071_),
    .C(_04098_),
    .Y(_03425_)
  );
  OAI21X1 _10680_ (
    .A(_03727_),
    .B(_04071_),
    .C(_04149_),
    .Y(_03390_)
  );
  OAI21X1 _10681_ (
    .A(_03728_),
    .B(_04071_),
    .C(_04150_),
    .Y(_03391_)
  );
  NAND2X1 _10682_ (
    .A(frontend_0.inst_jmp_bin_2_ ),
    .B(_04070_),
    .Y(_04158_)
  );
  OAI21X1 _10683_ (
    .A(_03706_),
    .B(_04070_),
    .C(_04158_),
    .Y(_03392_)
  );
  NAND2X1 _10684_ (
    .A(execution_unit_0.alu_0.inst_so_0_ ),
    .B(_04070_),
    .Y(_04159_)
  );
  AOI21X1 _10685_ (
    .A(_04145_),
    .B(_04159_),
    .C(_04108_),
    .Y(_03410_)
  );
  NAND2X1 _10686_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(_04070_),
    .Y(_04160_)
  );
  NAND3X1 _10687_ (
    .A(_03670_),
    .B(_03808_),
    .C(_04071_),
    .Y(_04161_)
  );
  OAI21X1 _10688_ (
    .A(_03672_),
    .B(_04161_),
    .C(_04160_),
    .Y(_03411_)
  );
  NAND2X1 _10689_ (
    .A(execution_unit_0.alu_0.inst_so_3_ ),
    .B(_04070_),
    .Y(_04162_)
  );
  OAI21X1 _10690_ (
    .A(_03774_),
    .B(_04147_),
    .C(_04162_),
    .Y(_03412_)
  );
  NAND2X1 _10691_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .B(_04070_),
    .Y(_04163_)
  );
  OAI21X1 _10692_ (
    .A(_03797_),
    .B(_04145_),
    .C(_04163_),
    .Y(_03413_)
  );
  NAND3X1 _10693_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(_03671_),
    .C(dbg_0.fe_mdb_in_7_ ),
    .Y(_04164_)
  );
  NAND2X1 _10694_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B(_04070_),
    .Y(_04165_)
  );
  OAI21X1 _10695_ (
    .A(_04155_),
    .B(_04164_),
    .C(_04165_),
    .Y(_03414_)
  );
  NAND2X1 _10696_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_04070_),
    .Y(_04166_)
  );
  OAI21X1 _10697_ (
    .A(_03798_),
    .B(_04070_),
    .C(_04166_),
    .Y(_03415_)
  );
  NOR2X1 _10698_ (
    .A(execution_unit_0.alu_0.inst_so_7_ ),
    .B(_04071_),
    .Y(_04167_)
  );
  AOI21X1 _10699_ (
    .A(_03775_),
    .B(_04071_),
    .C(_04167_),
    .Y(_03416_)
  );
  MUX2X1 _10700_ (
    .A(execution_unit_0.inst_dext_0_ ),
    .B(dbg_0.fe_mdb_in_0_ ),
    .S(_03910_),
    .Y(_04168_)
  );
  INVX1 _10701_ (
    .A(_04168_),
    .Y(_03373_)
  );
  NAND2X1 _10702_ (
    .A(execution_unit_0.inst_dext_1_ ),
    .B(_03910_),
    .Y(_04169_)
  );
  NOR2X1 _10703_ (
    .A(frontend_0.i_state_0_ ),
    .B(_03436_),
    .Y(_04170_)
  );
  OAI21X1 _10704_ (
    .A(_03873_),
    .B(_03876_),
    .C(_04170_),
    .Y(_04171_)
  );
  NAND3X1 _10705_ (
    .A(_03872_),
    .B(_03873_),
    .C(_04170_),
    .Y(_04172_)
  );
  OAI21X1 _10706_ (
    .A(_03881_),
    .B(_04172_),
    .C(frontend_0.i_state_5_ ),
    .Y(_04173_)
  );
  OAI21X1 _10707_ (
    .A(execution_unit_0.inst_as_4_ ),
    .B(_04173_),
    .C(_03685_),
    .Y(_03439_)
  );
  AOI22X1 _10708_ (
    .A(frontend_0.i_state_5_ ),
    .B(execution_unit_0.inst_as_4_ ),
    .C(_03439_),
    .D(execution_unit_0.UNUSED_inst_ad_symb ),
    .Y(_03440_)
  );
  OR2X1 _10709_ (
    .A(dbg_0.fe_mdb_in_1_ ),
    .B(_03440_),
    .Y(_03441_)
  );
  XNOR2X1 _10710_ (
    .A(_03677_),
    .B(_03440_),
    .Y(_03442_)
  );
  OAI21X1 _10711_ (
    .A(_03910_),
    .B(_03442_),
    .C(_04169_),
    .Y(_03380_)
  );
  NAND2X1 _10712_ (
    .A(execution_unit_0.inst_dext_2_ ),
    .B(_03910_),
    .Y(_03443_)
  );
  NOR2X1 _10713_ (
    .A(dbg_0.fe_mdb_in_2_ ),
    .B(_03441_),
    .Y(_03444_)
  );
  XNOR2X1 _10714_ (
    .A(_03678_),
    .B(_03441_),
    .Y(_03445_)
  );
  OAI21X1 _10715_ (
    .A(_03910_),
    .B(_03445_),
    .C(_03443_),
    .Y(_03381_)
  );
  OAI21X1 _10716_ (
    .A(dbg_0.fe_mdb_in_2_ ),
    .B(_03441_),
    .C(dbg_0.fe_mdb_in_3_ ),
    .Y(_03446_)
  );
  NAND2X1 _10717_ (
    .A(_03679_),
    .B(_03444_),
    .Y(_03447_)
  );
  AND2X1 _10718_ (
    .A(_03446_),
    .B(_03447_),
    .Y(_03448_)
  );
  NAND2X1 _10719_ (
    .A(execution_unit_0.inst_dext_3_ ),
    .B(_03910_),
    .Y(_03449_)
  );
  OAI21X1 _10720_ (
    .A(_03910_),
    .B(_03448_),
    .C(_03449_),
    .Y(_03382_)
  );
  NAND2X1 _10721_ (
    .A(execution_unit_0.inst_dext_4_ ),
    .B(_03910_),
    .Y(_03450_)
  );
  XNOR2X1 _10722_ (
    .A(_03675_),
    .B(_03447_),
    .Y(_03451_)
  );
  OAI21X1 _10723_ (
    .A(_03910_),
    .B(_03451_),
    .C(_03450_),
    .Y(_03383_)
  );
  OAI21X1 _10724_ (
    .A(dbg_0.fe_mdb_in_4_ ),
    .B(_03447_),
    .C(dbg_0.fe_mdb_in_5_ ),
    .Y(_03452_)
  );
  NAND3X1 _10725_ (
    .A(_03679_),
    .B(_04126_),
    .C(_03444_),
    .Y(_03453_)
  );
  AND2X1 _10726_ (
    .A(_03452_),
    .B(_03453_),
    .Y(_03454_)
  );
  NAND2X1 _10727_ (
    .A(execution_unit_0.inst_dext_5_ ),
    .B(_03910_),
    .Y(_03455_)
  );
  OAI21X1 _10728_ (
    .A(_03910_),
    .B(_03454_),
    .C(_03455_),
    .Y(_03384_)
  );
  NAND2X1 _10729_ (
    .A(execution_unit_0.inst_dext_6_ ),
    .B(_03910_),
    .Y(_03456_)
  );
  NOR2X1 _10730_ (
    .A(dbg_0.fe_mdb_in_6_ ),
    .B(_03453_),
    .Y(_03457_)
  );
  XNOR2X1 _10731_ (
    .A(_03698_),
    .B(_03453_),
    .Y(_03458_)
  );
  OAI21X1 _10732_ (
    .A(_03910_),
    .B(_03458_),
    .C(_03456_),
    .Y(_03385_)
  );
  OAI21X1 _10733_ (
    .A(dbg_0.fe_mdb_in_6_ ),
    .B(_03453_),
    .C(dbg_0.fe_mdb_in_7_ ),
    .Y(_03459_)
  );
  NAND2X1 _10734_ (
    .A(_03672_),
    .B(_03457_),
    .Y(_03460_)
  );
  AND2X1 _10735_ (
    .A(_03459_),
    .B(_03460_),
    .Y(_03461_)
  );
  NAND2X1 _10736_ (
    .A(execution_unit_0.inst_dext_7_ ),
    .B(_03910_),
    .Y(_03462_)
  );
  OAI21X1 _10737_ (
    .A(_03910_),
    .B(_03461_),
    .C(_03462_),
    .Y(_03386_)
  );
  NAND2X1 _10738_ (
    .A(execution_unit_0.inst_dext_8_ ),
    .B(_03910_),
    .Y(_03463_)
  );
  NAND3X1 _10739_ (
    .A(_03671_),
    .B(_03672_),
    .C(_03457_),
    .Y(_03464_)
  );
  XNOR2X1 _10740_ (
    .A(_03671_),
    .B(_03460_),
    .Y(_03465_)
  );
  OAI21X1 _10741_ (
    .A(_03910_),
    .B(_03465_),
    .C(_03463_),
    .Y(_03387_)
  );
  OAI21X1 _10742_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(_03460_),
    .C(dbg_0.fe_mdb_in_9_ ),
    .Y(_03466_)
  );
  OR2X1 _10743_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(_03464_),
    .Y(_03467_)
  );
  AND2X1 _10744_ (
    .A(_03466_),
    .B(_03467_),
    .Y(_03468_)
  );
  NAND2X1 _10745_ (
    .A(execution_unit_0.inst_dext_9_ ),
    .B(_03910_),
    .Y(_03469_)
  );
  OAI21X1 _10746_ (
    .A(_03910_),
    .B(_03468_),
    .C(_03469_),
    .Y(_03388_)
  );
  NAND2X1 _10747_ (
    .A(execution_unit_0.inst_dext_10_ ),
    .B(_03910_),
    .Y(_03470_)
  );
  NOR2X1 _10748_ (
    .A(dbg_0.fe_mdb_in_10_ ),
    .B(_03467_),
    .Y(_03471_)
  );
  XOR2X1 _10749_ (
    .A(dbg_0.fe_mdb_in_10_ ),
    .B(_03467_),
    .Y(_03472_)
  );
  OAI21X1 _10750_ (
    .A(_03910_),
    .B(_03472_),
    .C(_03470_),
    .Y(_03374_)
  );
  XNOR2X1 _10751_ (
    .A(dbg_0.fe_mdb_in_11_ ),
    .B(_03471_),
    .Y(_03473_)
  );
  NAND2X1 _10752_ (
    .A(execution_unit_0.inst_dext_11_ ),
    .B(_03910_),
    .Y(_03474_)
  );
  OAI21X1 _10753_ (
    .A(_03910_),
    .B(_03473_),
    .C(_03474_),
    .Y(_03375_)
  );
  NAND2X1 _10754_ (
    .A(execution_unit_0.inst_dext_12_ ),
    .B(_03910_),
    .Y(_03475_)
  );
  NOR2X1 _10755_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(dbg_0.fe_mdb_in_6_ ),
    .Y(_03476_)
  );
  NAND3X1 _10756_ (
    .A(_03785_),
    .B(_04106_),
    .C(_03476_),
    .Y(_03477_)
  );
  NOR2X1 _10757_ (
    .A(_03453_),
    .B(_03477_),
    .Y(_03478_)
  );
  OAI21X1 _10758_ (
    .A(_03453_),
    .B(_03477_),
    .C(dbg_0.fe_mdb_in_12_ ),
    .Y(_03479_)
  );
  NAND2X1 _10759_ (
    .A(_03706_),
    .B(_03478_),
    .Y(_03480_)
  );
  AND2X1 _10760_ (
    .A(_03479_),
    .B(_03480_),
    .Y(_03481_)
  );
  OAI21X1 _10761_ (
    .A(_03910_),
    .B(_03481_),
    .C(_03475_),
    .Y(_03376_)
  );
  OR2X1 _10762_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(_03480_),
    .Y(_03482_)
  );
  XNOR2X1 _10763_ (
    .A(_03673_),
    .B(_03480_),
    .Y(_03483_)
  );
  NAND2X1 _10764_ (
    .A(execution_unit_0.inst_dext_13_ ),
    .B(_03910_),
    .Y(_03484_)
  );
  OAI21X1 _10765_ (
    .A(_03910_),
    .B(_03483_),
    .C(_03484_),
    .Y(_03377_)
  );
  NAND2X1 _10766_ (
    .A(execution_unit_0.inst_dext_14_ ),
    .B(_03910_),
    .Y(_03485_)
  );
  NOR2X1 _10767_ (
    .A(dbg_0.fe_mdb_in_14_ ),
    .B(_03482_),
    .Y(_03486_)
  );
  XNOR2X1 _10768_ (
    .A(_03674_),
    .B(_03482_),
    .Y(_03487_)
  );
  OAI21X1 _10769_ (
    .A(_03910_),
    .B(_03487_),
    .C(_03485_),
    .Y(_03378_)
  );
  XNOR2X1 _10770_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(_03486_),
    .Y(_03488_)
  );
  NAND2X1 _10771_ (
    .A(execution_unit_0.inst_dext_15_ ),
    .B(_03910_),
    .Y(_03489_)
  );
  OAI21X1 _10772_ (
    .A(_03910_),
    .B(_03488_),
    .C(_03489_),
    .Y(_03379_)
  );
  NOR2X1 _10773_ (
    .A(_04070_),
    .B(_04139_),
    .Y(_03490_)
  );
  NAND2X1 _10774_ (
    .A(dbg_0.fe_mdb_in_4_ ),
    .B(_03490_),
    .Y(_03491_)
  );
  OAI21X1 _10775_ (
    .A(execution_unit_0.inst_sext_0_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03492_)
  );
  INVX1 _10776_ (
    .A(_03492_),
    .Y(_03493_)
  );
  OAI21X1 _10777_ (
    .A(dbg_0.fe_mdb_in_0_ ),
    .B(_03849_),
    .C(_03493_),
    .Y(_03494_)
  );
  OAI21X1 _10778_ (
    .A(_04141_),
    .B(_03494_),
    .C(_03491_),
    .Y(_03394_)
  );
  OAI21X1 _10779_ (
    .A(execution_unit_0.inst_sext_1_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03495_)
  );
  AOI21X1 _10780_ (
    .A(_03848_),
    .B(_03442_),
    .C(_03495_),
    .Y(_03496_)
  );
  AOI21X1 _10781_ (
    .A(dbg_0.fe_mdb_in_0_ ),
    .B(_04156_),
    .C(_03496_),
    .Y(_03497_)
  );
  NAND2X1 _10782_ (
    .A(dbg_0.fe_mdb_in_5_ ),
    .B(_03490_),
    .Y(_03498_)
  );
  OAI21X1 _10783_ (
    .A(_04141_),
    .B(_03497_),
    .C(_03498_),
    .Y(_03401_)
  );
  NOR2X1 _10784_ (
    .A(_03794_),
    .B(_04137_),
    .Y(_03499_)
  );
  NOR2X1 _10785_ (
    .A(_03782_),
    .B(_03815_),
    .Y(_03500_)
  );
  NOR2X1 _10786_ (
    .A(_03499_),
    .B(_03500_),
    .Y(_03501_)
  );
  OAI21X1 _10787_ (
    .A(execution_unit_0.inst_sext_2_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03502_)
  );
  AOI21X1 _10788_ (
    .A(_03848_),
    .B(_03445_),
    .C(_03502_),
    .Y(_03503_)
  );
  AOI21X1 _10789_ (
    .A(dbg_0.fe_mdb_in_1_ ),
    .B(_04156_),
    .C(_03503_),
    .Y(_03504_)
  );
  MUX2X1 _10790_ (
    .A(_03501_),
    .B(_03504_),
    .S(_04141_),
    .Y(_03402_)
  );
  OAI21X1 _10791_ (
    .A(execution_unit_0.inst_sext_3_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03505_)
  );
  AOI21X1 _10792_ (
    .A(_03848_),
    .B(_03448_),
    .C(_03505_),
    .Y(_03506_)
  );
  AOI21X1 _10793_ (
    .A(dbg_0.fe_mdb_in_2_ ),
    .B(_04156_),
    .C(_03506_),
    .Y(_03507_)
  );
  MUX2X1 _10794_ (
    .A(_03782_),
    .B(_03507_),
    .S(_04141_),
    .Y(_03403_)
  );
  OAI21X1 _10795_ (
    .A(execution_unit_0.inst_sext_4_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03508_)
  );
  AOI21X1 _10796_ (
    .A(_03848_),
    .B(_03451_),
    .C(_03508_),
    .Y(_03509_)
  );
  AOI21X1 _10797_ (
    .A(dbg_0.fe_mdb_in_3_ ),
    .B(_04156_),
    .C(_03509_),
    .Y(_03510_)
  );
  NAND2X1 _10798_ (
    .A(_04141_),
    .B(_03500_),
    .Y(_03511_)
  );
  OAI21X1 _10799_ (
    .A(_04141_),
    .B(_03510_),
    .C(_03511_),
    .Y(_03404_)
  );
  OAI21X1 _10800_ (
    .A(execution_unit_0.inst_sext_5_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03512_)
  );
  AOI21X1 _10801_ (
    .A(_03848_),
    .B(_03454_),
    .C(_03512_),
    .Y(_03513_)
  );
  AOI21X1 _10802_ (
    .A(dbg_0.fe_mdb_in_4_ ),
    .B(_04156_),
    .C(_03513_),
    .Y(_03514_)
  );
  OAI21X1 _10803_ (
    .A(_04141_),
    .B(_03514_),
    .C(_03511_),
    .Y(_03405_)
  );
  OAI21X1 _10804_ (
    .A(execution_unit_0.inst_sext_6_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03515_)
  );
  AOI21X1 _10805_ (
    .A(_03848_),
    .B(_03458_),
    .C(_03515_),
    .Y(_03516_)
  );
  AOI21X1 _10806_ (
    .A(dbg_0.fe_mdb_in_5_ ),
    .B(_04156_),
    .C(_03516_),
    .Y(_03517_)
  );
  OAI21X1 _10807_ (
    .A(_04141_),
    .B(_03517_),
    .C(_03511_),
    .Y(_03406_)
  );
  OAI21X1 _10808_ (
    .A(execution_unit_0.inst_sext_7_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03518_)
  );
  AOI21X1 _10809_ (
    .A(_03848_),
    .B(_03461_),
    .C(_03518_),
    .Y(_03519_)
  );
  AOI21X1 _10810_ (
    .A(dbg_0.fe_mdb_in_6_ ),
    .B(_04156_),
    .C(_03519_),
    .Y(_03520_)
  );
  OAI21X1 _10811_ (
    .A(_04141_),
    .B(_03520_),
    .C(_03511_),
    .Y(_03407_)
  );
  OAI21X1 _10812_ (
    .A(execution_unit_0.inst_sext_8_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03521_)
  );
  AOI21X1 _10813_ (
    .A(_03848_),
    .B(_03465_),
    .C(_03521_),
    .Y(_03522_)
  );
  AOI21X1 _10814_ (
    .A(dbg_0.fe_mdb_in_7_ ),
    .B(_04156_),
    .C(_03522_),
    .Y(_03523_)
  );
  OAI21X1 _10815_ (
    .A(_04141_),
    .B(_03523_),
    .C(_03511_),
    .Y(_03408_)
  );
  OAI21X1 _10816_ (
    .A(execution_unit_0.inst_sext_9_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03524_)
  );
  AOI21X1 _10817_ (
    .A(_03848_),
    .B(_03468_),
    .C(_03524_),
    .Y(_03525_)
  );
  AOI21X1 _10818_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(_04156_),
    .C(_03525_),
    .Y(_03526_)
  );
  OAI21X1 _10819_ (
    .A(_04141_),
    .B(_03526_),
    .C(_03511_),
    .Y(_03409_)
  );
  OAI21X1 _10820_ (
    .A(execution_unit_0.inst_sext_10_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03527_)
  );
  AOI21X1 _10821_ (
    .A(_03848_),
    .B(_03472_),
    .C(_03527_),
    .Y(_03528_)
  );
  NOR2X1 _10822_ (
    .A(_03670_),
    .B(_04157_),
    .Y(_03529_)
  );
  NOR2X1 _10823_ (
    .A(_03528_),
    .B(_03529_),
    .Y(_03530_)
  );
  OAI21X1 _10824_ (
    .A(_04141_),
    .B(_03530_),
    .C(_03511_),
    .Y(_03395_)
  );
  OAI21X1 _10825_ (
    .A(execution_unit_0.inst_sext_11_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03531_)
  );
  AOI21X1 _10826_ (
    .A(_03848_),
    .B(_03473_),
    .C(_03531_),
    .Y(_03532_)
  );
  NOR2X1 _10827_ (
    .A(_03529_),
    .B(_03532_),
    .Y(_03533_)
  );
  OAI21X1 _10828_ (
    .A(_04141_),
    .B(_03533_),
    .C(_03511_),
    .Y(_03396_)
  );
  OAI21X1 _10829_ (
    .A(execution_unit_0.inst_sext_12_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03534_)
  );
  AOI21X1 _10830_ (
    .A(_03848_),
    .B(_03481_),
    .C(_03534_),
    .Y(_03535_)
  );
  NOR2X1 _10831_ (
    .A(_03529_),
    .B(_03535_),
    .Y(_03536_)
  );
  OAI21X1 _10832_ (
    .A(_04141_),
    .B(_03536_),
    .C(_03511_),
    .Y(_03397_)
  );
  OAI21X1 _10833_ (
    .A(execution_unit_0.inst_sext_13_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03537_)
  );
  AOI21X1 _10834_ (
    .A(_03848_),
    .B(_03483_),
    .C(_03537_),
    .Y(_03538_)
  );
  NOR2X1 _10835_ (
    .A(_03529_),
    .B(_03538_),
    .Y(_03539_)
  );
  OAI21X1 _10836_ (
    .A(_04141_),
    .B(_03539_),
    .C(_03511_),
    .Y(_03398_)
  );
  OAI21X1 _10837_ (
    .A(execution_unit_0.inst_sext_14_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03540_)
  );
  AOI21X1 _10838_ (
    .A(_03848_),
    .B(_03487_),
    .C(_03540_),
    .Y(_03541_)
  );
  NOR2X1 _10839_ (
    .A(_03529_),
    .B(_03541_),
    .Y(_03542_)
  );
  OAI21X1 _10840_ (
    .A(_04141_),
    .B(_03542_),
    .C(_03511_),
    .Y(_03399_)
  );
  OAI21X1 _10841_ (
    .A(execution_unit_0.inst_sext_15_ ),
    .B(_03848_),
    .C(_04157_),
    .Y(_03543_)
  );
  AOI21X1 _10842_ (
    .A(_03848_),
    .B(_03488_),
    .C(_03543_),
    .Y(_03544_)
  );
  NOR2X1 _10843_ (
    .A(_03529_),
    .B(_03544_),
    .Y(_03545_)
  );
  OAI21X1 _10844_ (
    .A(_04141_),
    .B(_03545_),
    .C(_03511_),
    .Y(_03400_)
  );
  NAND2X1 _10845_ (
    .A(_03666_),
    .B(_03750_),
    .Y(_03546_)
  );
  OR2X1 _10846_ (
    .A(irq_11_),
    .B(_03546_),
    .Y(_03547_)
  );
  NAND2X1 _10847_ (
    .A(irq_9_),
    .B(_03752_),
    .Y(_03548_)
  );
  OAI22X1 _10848_ (
    .A(1'h0),
    .B(_03750_),
    .C(_03547_),
    .D(_03548_),
    .Y(_03549_)
  );
  AOI21X1 _10849_ (
    .A(irq_12_),
    .B(_03661_),
    .C(1'h0),
    .Y(_03550_)
  );
  OAI21X1 _10850_ (
    .A(_03752_),
    .B(_03547_),
    .C(_03550_),
    .Y(_03551_)
  );
  AOI21X1 _10851_ (
    .A(_03752_),
    .B(_03753_),
    .C(_03546_),
    .Y(_03552_)
  );
  NOR2X1 _10852_ (
    .A(_03549_),
    .B(_03552_),
    .Y(_03553_)
  );
  NAND2X1 _10853_ (
    .A(irq_8_),
    .B(_03553_),
    .Y(_03554_)
  );
  NOR2X1 _10854_ (
    .A(_03551_),
    .B(_03554_),
    .Y(_03555_)
  );
  OR2X1 _10855_ (
    .A(_03549_),
    .B(_03555_),
    .Y(_03556_)
  );
  INVX1 _10856_ (
    .A(_03556_),
    .Y(_03557_)
  );
  AOI21X1 _10857_ (
    .A(irq_8_),
    .B(_03553_),
    .C(_03551_),
    .Y(_03558_)
  );
  NAND3X1 _10858_ (
    .A(irq_6_),
    .B(_03662_),
    .C(_03553_),
    .Y(_03559_)
  );
  AND2X1 _10859_ (
    .A(_03558_),
    .B(_03559_),
    .Y(_03560_)
  );
  INVX1 _10860_ (
    .A(_03560_),
    .Y(_03561_)
  );
  NOR2X1 _10861_ (
    .A(_03552_),
    .B(_03561_),
    .Y(_03562_)
  );
  NAND2X1 _10862_ (
    .A(irq_4_),
    .B(_03562_),
    .Y(_03563_)
  );
  NAND2X1 _10863_ (
    .A(irq_5_),
    .B(_03553_),
    .Y(_03564_)
  );
  NOR2X1 _10864_ (
    .A(_03555_),
    .B(_03564_),
    .Y(_03565_)
  );
  NAND2X1 _10865_ (
    .A(_03560_),
    .B(_03565_),
    .Y(_03566_)
  );
  NOR2X1 _10866_ (
    .A(_03556_),
    .B(_03563_),
    .Y(_03567_)
  );
  AND2X1 _10867_ (
    .A(_03553_),
    .B(_03558_),
    .Y(_03568_)
  );
  OAI21X1 _10868_ (
    .A(irq_6_),
    .B(irq_7_),
    .C(_03568_),
    .Y(_03569_)
  );
  NAND2X1 _10869_ (
    .A(_03566_),
    .B(_03569_),
    .Y(_03570_)
  );
  NAND3X1 _10870_ (
    .A(_03566_),
    .B(_03567_),
    .C(_03569_),
    .Y(_03571_)
  );
  NAND3X1 _10871_ (
    .A(_03560_),
    .B(_03565_),
    .C(_03569_),
    .Y(_03572_)
  );
  NAND3X1 _10872_ (
    .A(_03557_),
    .B(_03571_),
    .C(_03572_),
    .Y(_03573_)
  );
  NOR2X1 _10873_ (
    .A(_03567_),
    .B(_03570_),
    .Y(_03574_)
  );
  NAND2X1 _10874_ (
    .A(_03562_),
    .B(_03574_),
    .Y(_03575_)
  );
  NOR2X1 _10875_ (
    .A(_03573_),
    .B(_03575_),
    .Y(_03576_)
  );
  NAND3X1 _10876_ (
    .A(irq_2_),
    .B(_03663_),
    .C(_03576_),
    .Y(_03577_)
  );
  NAND3X1 _10877_ (
    .A(_03560_),
    .B(_03571_),
    .C(_03577_),
    .Y(_03578_)
  );
  NOR2X1 _10878_ (
    .A(_03767_),
    .B(_03578_),
    .Y(_03579_)
  );
  NAND2X1 _10879_ (
    .A(irq_3_),
    .B(_03576_),
    .Y(_03580_)
  );
  NOR2X1 _10880_ (
    .A(_03552_),
    .B(_03555_),
    .Y(_03581_)
  );
  NAND3X1 _10881_ (
    .A(_03577_),
    .B(_03580_),
    .C(_03581_),
    .Y(_03582_)
  );
  NOR2X1 _10882_ (
    .A(_03573_),
    .B(_03582_),
    .Y(_03583_)
  );
  NAND3X1 _10883_ (
    .A(_03574_),
    .B(_03577_),
    .C(_03580_),
    .Y(_03584_)
  );
  NOR2X1 _10884_ (
    .A(_03578_),
    .B(_03584_),
    .Y(_03585_)
  );
  AND2X1 _10885_ (
    .A(_03664_),
    .B(_03583_),
    .Y(_03586_)
  );
  NAND3X1 _10886_ (
    .A(irq_0_),
    .B(_03585_),
    .C(_03586_),
    .Y(_03587_)
  );
  NAND3X1 _10887_ (
    .A(irq_1_),
    .B(_03583_),
    .C(_03585_),
    .Y(_03588_)
  );
  NAND2X1 _10888_ (
    .A(_03579_),
    .B(_03587_),
    .Y(_03589_)
  );
  OAI21X1 _10889_ (
    .A(_03690_),
    .B(_03766_),
    .C(_03589_),
    .Y(_03426_)
  );
  NAND3X1 _10890_ (
    .A(_03766_),
    .B(_03587_),
    .C(_03588_),
    .Y(_03590_)
  );
  OAI22X1 _10891_ (
    .A(_03692_),
    .B(_03766_),
    .C(_03573_),
    .D(_03590_),
    .Y(_03427_)
  );
  OAI22X1 _10892_ (
    .A(_03694_),
    .B(_03766_),
    .C(_03582_),
    .D(_03590_),
    .Y(_03428_)
  );
  OAI21X1 _10893_ (
    .A(_03749_),
    .B(_03765_),
    .C(frontend_0.irq_addr_4_ ),
    .Y(_03591_)
  );
  OAI21X1 _10894_ (
    .A(_03584_),
    .B(_03590_),
    .C(_03591_),
    .Y(_03429_)
  );
  OR2X1 _10895_ (
    .A(frontend_0.irq_addr_5_ ),
    .B(_03766_),
    .Y(_03430_)
  );
  OAI21X1 _10896_ (
    .A(_03749_),
    .B(_03765_),
    .C(_03699_),
    .Y(_03431_)
  );
  NOR2X1 _10897_ (
    .A(_03729_),
    .B(exec_done),
    .Y(_03389_)
  );
  OAI21X1 _10898_ (
    .A(_03436_),
    .B(_03432_),
    .C(_03762_),
    .Y(_03592_)
  );
  NOR2X1 _10899_ (
    .A(_03874_),
    .B(_03592_),
    .Y(_03593_)
  );
  NAND2X1 _10900_ (
    .A(_04171_),
    .B(_03593_),
    .Y(_03594_)
  );
  INVX1 _10901_ (
    .A(_03594_),
    .Y(_03340_)
  );
  AND2X1 _10902_ (
    .A(frontend_0.irq_addr_5_ ),
    .B(frontend_0.irq_addr_6_ ),
    .Y(_03595_)
  );
  NAND2X1 _10903_ (
    .A(frontend_0.irq_addr_5_ ),
    .B(frontend_0.irq_addr_6_ ),
    .Y(_03596_)
  );
  NOR2X1 _10904_ (
    .A(_03690_),
    .B(frontend_0.irq_addr_2_ ),
    .Y(_03597_)
  );
  NAND2X1 _10905_ (
    .A(frontend_0.irq_addr_1_ ),
    .B(_03692_),
    .Y(_03598_)
  );
  AND2X1 _10906_ (
    .A(frontend_0.irq_addr_3_ ),
    .B(frontend_0.irq_addr_4_ ),
    .Y(_03599_)
  );
  NAND2X1 _10907_ (
    .A(_03597_),
    .B(_03599_),
    .Y(_03600_)
  );
  NAND2X1 _10908_ (
    .A(frontend_0.irq_addr_1_ ),
    .B(frontend_0.irq_addr_2_ ),
    .Y(_03601_)
  );
  INVX1 _10909_ (
    .A(_03601_),
    .Y(_03602_)
  );
  NAND2X1 _10910_ (
    .A(_03694_),
    .B(frontend_0.irq_addr_4_ ),
    .Y(_03603_)
  );
  OAI21X1 _10911_ (
    .A(_03601_),
    .B(_03603_),
    .C(_03600_),
    .Y(_03604_)
  );
  NAND2X1 _10912_ (
    .A(_03595_),
    .B(_03604_),
    .Y(_03605_)
  );
  NAND3X1 _10913_ (
    .A(_03595_),
    .B(_03598_),
    .C(_03599_),
    .Y(_03606_)
  );
  NOR2X1 _10914_ (
    .A(_03596_),
    .B(_03603_),
    .Y(_03607_)
  );
  OR2X1 _10915_ (
    .A(_03596_),
    .B(_03603_),
    .Y(_03608_)
  );
  NOR2X1 _10916_ (
    .A(frontend_0.irq_addr_1_ ),
    .B(frontend_0.irq_addr_2_ ),
    .Y(_03609_)
  );
  INVX1 _10917_ (
    .A(_03609_),
    .Y(_03610_)
  );
  NOR2X1 _10918_ (
    .A(frontend_0.irq_addr_1_ ),
    .B(_03692_),
    .Y(_03611_)
  );
  NAND2X1 _10919_ (
    .A(_03690_),
    .B(frontend_0.irq_addr_2_ ),
    .Y(_03612_)
  );
  OAI21X1 _10920_ (
    .A(_03597_),
    .B(_03611_),
    .C(_03607_),
    .Y(_03613_)
  );
  NAND3X1 _10921_ (
    .A(_03605_),
    .B(_03606_),
    .C(_03613_),
    .Y(_03614_)
  );
  OR2X1 _10922_ (
    .A(_03603_),
    .B(_03610_),
    .Y(_03615_)
  );
  NOR2X1 _10923_ (
    .A(_03694_),
    .B(frontend_0.irq_addr_4_ ),
    .Y(_03616_)
  );
  OAI21X1 _10924_ (
    .A(frontend_0.irq_addr_1_ ),
    .B(frontend_0.irq_addr_2_ ),
    .C(_03616_),
    .Y(_03617_)
  );
  AOI21X1 _10925_ (
    .A(_03615_),
    .B(_03617_),
    .C(_03596_),
    .Y(_03618_)
  );
  OR2X1 _10926_ (
    .A(_03614_),
    .B(_03618_),
    .Y(_03619_)
  );
  NOR2X1 _10927_ (
    .A(frontend_0.irq_addr_3_ ),
    .B(frontend_0.irq_addr_4_ ),
    .Y(_03620_)
  );
  AOI22X1 _10928_ (
    .A(_03609_),
    .B(_03616_),
    .C(_03620_),
    .D(_03602_),
    .Y(_03621_)
  );
  NOR2X1 _10929_ (
    .A(_03699_),
    .B(_03954_),
    .Y(_03622_)
  );
  OR2X1 _10930_ (
    .A(_03699_),
    .B(_03954_),
    .Y(_03623_)
  );
  OAI21X1 _10931_ (
    .A(_03597_),
    .B(_03611_),
    .C(_03620_),
    .Y(_03624_)
  );
  AND2X1 _10932_ (
    .A(_03622_),
    .B(_03624_),
    .Y(_03625_)
  );
  OAI21X1 _10933_ (
    .A(_03596_),
    .B(_03621_),
    .C(_03625_),
    .Y(_03626_)
  );
  NOR2X1 _10934_ (
    .A(_03619_),
    .B(_03626_),
    .Y(_00083_)
  );
  OR2X1 _10935_ (
    .A(_03619_),
    .B(_03623_),
    .Y(_03627_)
  );
  INVX1 _10936_ (
    .A(_03627_),
    .Y(_03628_)
  );
  NAND2X1 _10937_ (
    .A(_03621_),
    .B(_03628_),
    .Y(_03629_)
  );
  AOI21X1 _10938_ (
    .A(_03690_),
    .B(_03620_),
    .C(_03629_),
    .Y(_00088_)
  );
  NAND2X1 _10939_ (
    .A(_03595_),
    .B(_03620_),
    .Y(_03630_)
  );
  NOR2X1 _10940_ (
    .A(frontend_0.irq_addr_2_ ),
    .B(_03630_),
    .Y(_03631_)
  );
  NOR2X1 _10941_ (
    .A(_03629_),
    .B(_03631_),
    .Y(_00089_)
  );
  AOI22X1 _10942_ (
    .A(_03609_),
    .B(_03616_),
    .C(_03620_),
    .D(_03611_),
    .Y(_03632_)
  );
  OAI21X1 _10943_ (
    .A(frontend_0.irq_addr_2_ ),
    .B(_03630_),
    .C(_03632_),
    .Y(_03633_)
  );
  NOR2X1 _10944_ (
    .A(_03627_),
    .B(_03633_),
    .Y(_00090_)
  );
  NOR2X1 _10945_ (
    .A(_03620_),
    .B(_03627_),
    .Y(_00091_)
  );
  NAND3X1 _10946_ (
    .A(_03615_),
    .B(_03622_),
    .C(_03630_),
    .Y(_03634_)
  );
  OR2X1 _10947_ (
    .A(_03614_),
    .B(_03634_),
    .Y(_03635_)
  );
  AOI21X1 _10948_ (
    .A(_03598_),
    .B(_03616_),
    .C(_03635_),
    .Y(_00092_)
  );
  OAI21X1 _10949_ (
    .A(frontend_0.irq_addr_2_ ),
    .B(_03596_),
    .C(_03601_),
    .Y(_03636_)
  );
  AOI21X1 _10950_ (
    .A(_03616_),
    .B(_03636_),
    .C(_03635_),
    .Y(_00093_)
  );
  OAI21X1 _10951_ (
    .A(frontend_0.irq_addr_2_ ),
    .B(_03596_),
    .C(_03612_),
    .Y(_03637_)
  );
  AOI21X1 _10952_ (
    .A(_03616_),
    .B(_03637_),
    .C(_03635_),
    .Y(_00094_)
  );
  NAND3X1 _10953_ (
    .A(frontend_0.irq_addr_4_ ),
    .B(_03606_),
    .C(_03622_),
    .Y(_03638_)
  );
  INVX1 _10954_ (
    .A(_03638_),
    .Y(_03639_)
  );
  NOR2X1 _10955_ (
    .A(_03604_),
    .B(_03638_),
    .Y(_03640_)
  );
  AND2X1 _10956_ (
    .A(_03613_),
    .B(_03640_),
    .Y(_00095_)
  );
  OAI21X1 _10957_ (
    .A(frontend_0.irq_addr_1_ ),
    .B(_03608_),
    .C(_03640_),
    .Y(_03641_)
  );
  INVX1 _10958_ (
    .A(_03641_),
    .Y(_00096_)
  );
  OAI21X1 _10959_ (
    .A(frontend_0.irq_addr_2_ ),
    .B(_03608_),
    .C(_03639_),
    .Y(_03642_)
  );
  AOI21X1 _10960_ (
    .A(_03595_),
    .B(_03604_),
    .C(_03642_),
    .Y(_00084_)
  );
  OAI21X1 _10961_ (
    .A(_03603_),
    .B(_03612_),
    .C(_03600_),
    .Y(_03643_)
  );
  AOI21X1 _10962_ (
    .A(_03595_),
    .B(_03643_),
    .C(_03642_),
    .Y(_00085_)
  );
  NAND2X1 _10963_ (
    .A(_03599_),
    .B(_03622_),
    .Y(_03644_)
  );
  NOR2X1 _10964_ (
    .A(_03610_),
    .B(_03644_),
    .Y(_00086_)
  );
  NOR2X1 _10965_ (
    .A(_03600_),
    .B(_03623_),
    .Y(_00087_)
  );
  OR2X1 _10966_ (
    .A(frontend_0.pmem_busy ),
    .B(_03882_),
    .Y(_03645_)
  );
  AOI21X1 _10967_ (
    .A(cpu_halt_st),
    .B(_03761_),
    .C(_03645_),
    .Y(_03646_)
  );
  OAI21X1 _10968_ (
    .A(_03863_),
    .B(_03920_),
    .C(_03646_),
    .Y(fe_mb_en)
  );
  OR2X1 _10969_ (
    .A(_03714_),
    .B(frontend_0.inst_jmp_bin_2_ ),
    .Y(_03647_)
  );
  NAND2X1 _10970_ (
    .A(_03727_),
    .B(_03728_),
    .Y(_03648_)
  );
  NOR2X1 _10971_ (
    .A(_03647_),
    .B(_03648_),
    .Y(execution_unit_0.alu_0.inst_jmp_0_ )
  );
  NAND2X1 _10972_ (
    .A(frontend_0.inst_jmp_bin_0_ ),
    .B(_03728_),
    .Y(_03649_)
  );
  NOR2X1 _10973_ (
    .A(_03647_),
    .B(_03649_),
    .Y(execution_unit_0.alu_0.inst_jmp_1_ )
  );
  NAND2X1 _10974_ (
    .A(_03727_),
    .B(frontend_0.inst_jmp_bin_1_ ),
    .Y(_03650_)
  );
  NOR2X1 _10975_ (
    .A(_03647_),
    .B(_03650_),
    .Y(execution_unit_0.alu_0.inst_jmp_2_ )
  );
  NAND2X1 _10976_ (
    .A(frontend_0.inst_jmp_bin_0_ ),
    .B(frontend_0.inst_jmp_bin_1_ ),
    .Y(_03651_)
  );
  NOR2X1 _10977_ (
    .A(_03647_),
    .B(_03651_),
    .Y(execution_unit_0.alu_0.inst_jmp_3_ )
  );
  NAND2X1 _10978_ (
    .A(execution_unit_0.inst_type_1_ ),
    .B(frontend_0.inst_jmp_bin_2_ ),
    .Y(_03652_)
  );
  NOR2X1 _10979_ (
    .A(_03648_),
    .B(_03652_),
    .Y(execution_unit_0.alu_0.inst_jmp_4_ )
  );
  NOR2X1 _10980_ (
    .A(_03649_),
    .B(_03652_),
    .Y(execution_unit_0.alu_0.inst_jmp_5_ )
  );
  NOR2X1 _10981_ (
    .A(_03650_),
    .B(_03652_),
    .Y(execution_unit_0.alu_0.inst_jmp_6_ )
  );
  NAND2X1 _10982_ (
    .A(execution_unit_0.inst_type_0_ ),
    .B(_03837_),
    .Y(_03653_)
  );
  OAI21X1 _10983_ (
    .A(_03736_),
    .B(_03737_),
    .C(frontend_0.exec_src_wr ),
    .Y(_03654_)
  );
  OAI21X1 _10984_ (
    .A(_03744_),
    .B(_03654_),
    .C(_03653_),
    .Y(_03344_)
  );
  OAI21X1 _10985_ (
    .A(_03736_),
    .B(_03828_),
    .C(_03740_),
    .Y(_03342_)
  );
  NOR2X1 _10986_ (
    .A(dbg_0.fe_mdb_in_7_ ),
    .B(_04118_),
    .Y(_03655_)
  );
  AOI21X1 _10987_ (
    .A(_03806_),
    .B(_03655_),
    .C(_04091_),
    .Y(_03656_)
  );
  OAI21X1 _10988_ (
    .A(_04070_),
    .B(_03656_),
    .C(_03733_),
    .Y(_03343_)
  );
  DFFSR _10989_ (
    .CLK(dco_clk),
    .D(_03434_),
    .Q(frontend_0.i_state_0_ ),
    .R(1'h1),
    .S(_03438_)
  );
  DFFSR _10990_ (
    .CLK(dco_clk),
    .D(_03432_),
    .Q(frontend_0.i_state_1_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _10991_ (
    .CLK(dco_clk),
    .D(_03435_),
    .Q(frontend_0.i_state_2_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _10992_ (
    .CLK(dco_clk),
    .D(frontend_0.i_state_0_ ),
    .Q(frontend_0.i_state_3_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _10993_ (
    .CLK(dco_clk),
    .D(_03436_),
    .Q(frontend_0.i_state_4_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _10994_ (
    .CLK(dco_clk),
    .D(_03433_),
    .Q(frontend_0.i_state_5_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _10995_ (
    .CLK(dco_clk),
    .D(_03349_),
    .Q(execution_unit_0.alu_0.inst_alu_0_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _10996_ (
    .CLK(dco_clk),
    .D(_03351_),
    .Q(execution_unit_0.alu_0.inst_alu_1_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _10997_ (
    .CLK(dco_clk),
    .D(_03352_),
    .Q(execution_unit_0.alu_0.inst_alu_2_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _10998_ (
    .CLK(dco_clk),
    .D(_03353_),
    .Q(execution_unit_0.alu_0.inst_alu_3_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _10999_ (
    .CLK(dco_clk),
    .D(_03354_),
    .Q(execution_unit_0.alu_0.inst_alu_4_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11000_ (
    .CLK(dco_clk),
    .D(_03355_),
    .Q(execution_unit_0.alu_0.inst_alu_5_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11001_ (
    .CLK(dco_clk),
    .D(_03356_),
    .Q(execution_unit_0.alu_0.inst_alu_6_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11002_ (
    .CLK(dco_clk),
    .D(_03357_),
    .Q(execution_unit_0.alu_0.inst_alu_7_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11003_ (
    .CLK(dco_clk),
    .D(_03358_),
    .Q(execution_unit_0.alu_0.inst_alu_8_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11004_ (
    .CLK(dco_clk),
    .D(_03359_),
    .Q(execution_unit_0.alu_0.inst_alu_9_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11005_ (
    .CLK(dco_clk),
    .D(_03350_),
    .Q(execution_unit_0.alu_0.inst_alu_10_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11006_ (
    .CLK(dco_clk),
    .D(_03437_),
    .Q(execution_unit_0.alu_0.UNUSED_inst_alu ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11007_ (
    .CLK(dco_clk),
    .D(frontend_0.e_state_nxt_0_ ),
    .Q(e_state_0_),
    .R(1'h1),
    .S(_03438_)
  );
  DFFSR _11008_ (
    .CLK(dco_clk),
    .D(frontend_0.e_state_nxt_1_ ),
    .Q(e_state_1_),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11009_ (
    .CLK(dco_clk),
    .D(frontend_0.e_state_nxt_2_ ),
    .Q(e_state_2_),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11010_ (
    .CLK(dco_clk),
    .D(frontend_0.e_state_nxt_3_ ),
    .Q(e_state_3_),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11011_ (
    .CLK(dco_clk),
    .D(_03341_),
    .Q(frontend_0.exec_dext_rdy ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11012_ (
    .CLK(dco_clk),
    .D(_03344_),
    .Q(frontend_0.exec_src_wr ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11013_ (
    .CLK(dco_clk),
    .D(_03342_),
    .Q(frontend_0.exec_dst_wr ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11014_ (
    .CLK(dco_clk),
    .D(_03343_),
    .Q(frontend_0.exec_jmp ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11015_ (
    .CLK(dco_clk),
    .D(_03421_),
    .Q(frontend_0.inst_sz_0_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11016_ (
    .CLK(dco_clk),
    .D(_03422_),
    .Q(frontend_0.inst_sz_1_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11017_ (
    .CLK(dco_clk),
    .D(_03368_),
    .Q(execution_unit_0.alu_0.inst_bw ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11018_ (
    .CLK(dco_clk),
    .D(_03345_),
    .Q(execution_unit_0.inst_ad_0_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11019_ (
    .CLK(dco_clk),
    .D(_03346_),
    .Q(execution_unit_0.UNUSED_inst_ad_idx ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11020_ (
    .CLK(dco_clk),
    .D(_03347_),
    .Q(execution_unit_0.UNUSED_inst_ad_symb ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11021_ (
    .CLK(dco_clk),
    .D(_03348_),
    .Q(execution_unit_0.inst_ad_6_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11022_ (
    .CLK(dco_clk),
    .D(_03360_),
    .Q(execution_unit_0.inst_as_0_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11023_ (
    .CLK(dco_clk),
    .D(_03361_),
    .Q(execution_unit_0.inst_as_1_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11024_ (
    .CLK(dco_clk),
    .D(_03362_),
    .Q(execution_unit_0.inst_as_2_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11025_ (
    .CLK(dco_clk),
    .D(_03363_),
    .Q(execution_unit_0.inst_as_3_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11026_ (
    .CLK(dco_clk),
    .D(_03364_),
    .Q(execution_unit_0.inst_as_4_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11027_ (
    .CLK(dco_clk),
    .D(_03365_),
    .Q(execution_unit_0.inst_as_5_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11028_ (
    .CLK(dco_clk),
    .D(_03366_),
    .Q(execution_unit_0.inst_as_6_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11029_ (
    .CLK(dco_clk),
    .D(_03367_),
    .Q(execution_unit_0.inst_as_7_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11030_ (
    .CLK(dco_clk),
    .D(_03417_),
    .Q(frontend_0.inst_src_bin_0_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11031_ (
    .CLK(dco_clk),
    .D(_03418_),
    .Q(frontend_0.inst_src_bin_1_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11032_ (
    .CLK(dco_clk),
    .D(_03419_),
    .Q(frontend_0.inst_src_bin_2_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11033_ (
    .CLK(dco_clk),
    .D(_03420_),
    .Q(frontend_0.inst_src_bin_3_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11034_ (
    .CLK(dco_clk),
    .D(_03369_),
    .Q(frontend_0.inst_dest_bin_0_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11035_ (
    .CLK(dco_clk),
    .D(_03370_),
    .Q(frontend_0.inst_dest_bin_1_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11036_ (
    .CLK(dco_clk),
    .D(_03371_),
    .Q(frontend_0.inst_dest_bin_2_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11037_ (
    .CLK(dco_clk),
    .D(_03372_),
    .Q(frontend_0.inst_dest_bin_3_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11038_ (
    .CLK(dco_clk),
    .D(_03393_),
    .Q(execution_unit_0.inst_mov ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11039_ (
    .CLK(dco_clk),
    .D(_03390_),
    .Q(frontend_0.inst_jmp_bin_0_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11040_ (
    .CLK(dco_clk),
    .D(_03391_),
    .Q(frontend_0.inst_jmp_bin_1_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11041_ (
    .CLK(dco_clk),
    .D(_03392_),
    .Q(frontend_0.inst_jmp_bin_2_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11042_ (
    .CLK(dco_clk),
    .D(_03410_),
    .Q(execution_unit_0.alu_0.inst_so_0_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11043_ (
    .CLK(dco_clk),
    .D(_03411_),
    .Q(execution_unit_0.alu_0.inst_so_1_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11044_ (
    .CLK(dco_clk),
    .D(_03412_),
    .Q(execution_unit_0.alu_0.inst_so_3_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11045_ (
    .CLK(dco_clk),
    .D(_03413_),
    .Q(execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11046_ (
    .CLK(dco_clk),
    .D(_03414_),
    .Q(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11047_ (
    .CLK(dco_clk),
    .D(_03415_),
    .Q(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11048_ (
    .CLK(dco_clk),
    .D(_03416_),
    .Q(execution_unit_0.alu_0.inst_so_7_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11049_ (
    .CLK(dco_clk),
    .D(_03423_),
    .Q(execution_unit_0.inst_type_0_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11050_ (
    .CLK(dco_clk),
    .D(_03424_),
    .Q(execution_unit_0.inst_type_1_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11051_ (
    .CLK(dco_clk),
    .D(_03425_),
    .Q(execution_unit_0.inst_type_2_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11052_ (
    .CLK(dco_clk),
    .D(_03373_),
    .Q(execution_unit_0.inst_dext_0_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11053_ (
    .CLK(dco_clk),
    .D(_03380_),
    .Q(execution_unit_0.inst_dext_1_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11054_ (
    .CLK(dco_clk),
    .D(_03381_),
    .Q(execution_unit_0.inst_dext_2_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11055_ (
    .CLK(dco_clk),
    .D(_03382_),
    .Q(execution_unit_0.inst_dext_3_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11056_ (
    .CLK(dco_clk),
    .D(_03383_),
    .Q(execution_unit_0.inst_dext_4_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11057_ (
    .CLK(dco_clk),
    .D(_03384_),
    .Q(execution_unit_0.inst_dext_5_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11058_ (
    .CLK(dco_clk),
    .D(_03385_),
    .Q(execution_unit_0.inst_dext_6_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11059_ (
    .CLK(dco_clk),
    .D(_03386_),
    .Q(execution_unit_0.inst_dext_7_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11060_ (
    .CLK(dco_clk),
    .D(_03387_),
    .Q(execution_unit_0.inst_dext_8_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11061_ (
    .CLK(dco_clk),
    .D(_03388_),
    .Q(execution_unit_0.inst_dext_9_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11062_ (
    .CLK(dco_clk),
    .D(_03374_),
    .Q(execution_unit_0.inst_dext_10_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11063_ (
    .CLK(dco_clk),
    .D(_03375_),
    .Q(execution_unit_0.inst_dext_11_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11064_ (
    .CLK(dco_clk),
    .D(_03376_),
    .Q(execution_unit_0.inst_dext_12_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11065_ (
    .CLK(dco_clk),
    .D(_03377_),
    .Q(execution_unit_0.inst_dext_13_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11066_ (
    .CLK(dco_clk),
    .D(_03378_),
    .Q(execution_unit_0.inst_dext_14_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11067_ (
    .CLK(dco_clk),
    .D(_03379_),
    .Q(execution_unit_0.inst_dext_15_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11068_ (
    .CLK(dco_clk),
    .D(_03394_),
    .Q(execution_unit_0.inst_sext_0_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11069_ (
    .CLK(dco_clk),
    .D(_03401_),
    .Q(execution_unit_0.inst_sext_1_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11070_ (
    .CLK(dco_clk),
    .D(_03402_),
    .Q(execution_unit_0.inst_sext_2_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11071_ (
    .CLK(dco_clk),
    .D(_03403_),
    .Q(execution_unit_0.inst_sext_3_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11072_ (
    .CLK(dco_clk),
    .D(_03404_),
    .Q(execution_unit_0.inst_sext_4_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11073_ (
    .CLK(dco_clk),
    .D(_03405_),
    .Q(execution_unit_0.inst_sext_5_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11074_ (
    .CLK(dco_clk),
    .D(_03406_),
    .Q(execution_unit_0.inst_sext_6_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11075_ (
    .CLK(dco_clk),
    .D(_03407_),
    .Q(execution_unit_0.inst_sext_7_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11076_ (
    .CLK(dco_clk),
    .D(_03408_),
    .Q(execution_unit_0.inst_sext_8_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11077_ (
    .CLK(dco_clk),
    .D(_03409_),
    .Q(execution_unit_0.inst_sext_9_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11078_ (
    .CLK(dco_clk),
    .D(_03395_),
    .Q(execution_unit_0.inst_sext_10_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11079_ (
    .CLK(dco_clk),
    .D(_03396_),
    .Q(execution_unit_0.inst_sext_11_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11080_ (
    .CLK(dco_clk),
    .D(_03397_),
    .Q(execution_unit_0.inst_sext_12_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11081_ (
    .CLK(dco_clk),
    .D(_03398_),
    .Q(execution_unit_0.inst_sext_13_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11082_ (
    .CLK(dco_clk),
    .D(_03399_),
    .Q(execution_unit_0.inst_sext_14_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11083_ (
    .CLK(dco_clk),
    .D(_03400_),
    .Q(execution_unit_0.inst_sext_15_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11084_ (
    .CLK(dco_clk),
    .D(fe_pmem_wait),
    .Q(frontend_0.pmem_busy ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11085_ (
    .CLK(dco_clk),
    .D(UNUSED_fe_mab_0),
    .Q(dbg_0.UNUSED_pc_0_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11086_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_1_ ),
    .Q(dbg_0.UNUSED_pc_1_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11087_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_2_ ),
    .Q(dbg_0.UNUSED_pc_2_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11088_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_3_ ),
    .Q(dbg_0.UNUSED_pc_3_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11089_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_4_ ),
    .Q(dbg_0.UNUSED_pc_4_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11090_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_5_ ),
    .Q(dbg_0.UNUSED_pc_5_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11091_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_6_ ),
    .Q(dbg_0.UNUSED_pc_6_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11092_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_7_ ),
    .Q(dbg_0.UNUSED_pc_7_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11093_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_8_ ),
    .Q(dbg_0.UNUSED_pc_8_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11094_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_9_ ),
    .Q(dbg_0.UNUSED_pc_9_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11095_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_10_ ),
    .Q(dbg_0.UNUSED_pc_10_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11096_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_11_ ),
    .Q(dbg_0.UNUSED_pc_11_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11097_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_12_ ),
    .Q(dbg_0.UNUSED_pc_12_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11098_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_13_ ),
    .Q(dbg_0.UNUSED_pc_13_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11099_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_14_ ),
    .Q(dbg_0.UNUSED_pc_14_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11100_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_15_ ),
    .Q(dbg_0.UNUSED_pc_15_ ),
    .R(_03438_),
    .S(1'h1)
  );
  DFFSR _11101_ (
    .CLK(dco_clk),
    .D(_03426_),
    .Q(frontend_0.irq_addr_1_ ),
    .R(1'h1),
    .S(_03438_)
  );
  DFFSR _11102_ (
    .CLK(dco_clk),
    .D(_03427_),
    .Q(frontend_0.irq_addr_2_ ),
    .R(1'h1),
    .S(_03438_)
  );
  DFFSR _11103_ (
    .CLK(dco_clk),
    .D(_03428_),
    .Q(frontend_0.irq_addr_3_ ),
    .R(1'h1),
    .S(_03438_)
  );
  DFFSR _11104_ (
    .CLK(dco_clk),
    .D(_03429_),
    .Q(frontend_0.irq_addr_4_ ),
    .R(1'h1),
    .S(_03438_)
  );
  DFFSR _11105_ (
    .CLK(dco_clk),
    .D(_03430_),
    .Q(frontend_0.irq_addr_5_ ),
    .R(1'h1),
    .S(_03438_)
  );
  DFFSR _11106_ (
    .CLK(dco_clk),
    .D(_03431_),
    .Q(frontend_0.irq_addr_6_ ),
    .R(1'h1),
    .S(_03438_)
  );
  DFFSR _11107_ (
    .CLK(dco_clk),
    .D(_03389_),
    .Q(execution_unit_0.inst_irq_rst ),
    .R(1'h1),
    .S(_03438_)
  );
  DFFSR _11108_ (
    .CLK(dco_clk),
    .D(_03340_),
    .Q(cpu_halt_st),
    .R(_03438_),
    .S(1'h1)
  );
  INVX1 _11109_ (
    .A(dbg_0.UNUSED_eu_mb_wr_1_ ),
    .Y(_04192_)
  );
  INVX1 _11110_ (
    .A(dbg_0.dbg_mem_wr_1_ ),
    .Y(_04193_)
  );
  INVX1 _11111_ (
    .A(dbg_0.dbg_mem_addr_15_ ),
    .Y(_04194_)
  );
  INVX1 _11112_ (
    .A(dbg_0.dbg_mem_addr_14_ ),
    .Y(_04195_)
  );
  INVX1 _11113_ (
    .A(dbg_0.dbg_mem_addr_13_ ),
    .Y(_04196_)
  );
  INVX1 _11114_ (
    .A(dbg_0.dbg_mem_addr_12_ ),
    .Y(_04197_)
  );
  INVX1 _11115_ (
    .A(dbg_0.dbg_mem_addr_11_ ),
    .Y(_04198_)
  );
  INVX1 _11116_ (
    .A(dbg_0.dbg_mem_addr_10_ ),
    .Y(_04199_)
  );
  INVX1 _11117_ (
    .A(dbg_0.dbg_mem_addr_9_ ),
    .Y(_04200_)
  );
  INVX1 _11118_ (
    .A(dbg_0.dbg_mem_addr_8_ ),
    .Y(_04201_)
  );
  INVX1 _11119_ (
    .A(dbg_0.dbg_mem_addr_7_ ),
    .Y(_04202_)
  );
  INVX1 _11120_ (
    .A(dbg_0.dbg_mem_addr_6_ ),
    .Y(_04203_)
  );
  INVX1 _11121_ (
    .A(dbg_0.dbg_mem_addr_5_ ),
    .Y(_04204_)
  );
  INVX1 _11122_ (
    .A(dbg_0.dbg_mem_addr_4_ ),
    .Y(_04205_)
  );
  INVX1 _11123_ (
    .A(dbg_0.dbg_mem_addr_3_ ),
    .Y(_04206_)
  );
  INVX1 _11124_ (
    .A(dbg_0.dbg_mem_addr_2_ ),
    .Y(_04207_)
  );
  INVX1 _11125_ (
    .A(dbg_0.dbg_mem_addr_1_ ),
    .Y(_04208_)
  );
  INVX1 _11126_ (
    .A(dbg_0.UNUSED_eu_mb_en ),
    .Y(_04209_)
  );
  INVX1 _11127_ (
    .A(dbg_0.UNUSED_eu_mab_13_ ),
    .Y(_04210_)
  );
  INVX1 _11128_ (
    .A(dbg_0.UNUSED_eu_mab_12_ ),
    .Y(_04211_)
  );
  INVX1 _11129_ (
    .A(dbg_0.UNUSED_eu_mab_11_ ),
    .Y(_04212_)
  );
  INVX1 _11130_ (
    .A(dbg_0.UNUSED_eu_mab_10_ ),
    .Y(_04213_)
  );
  INVX1 _11131_ (
    .A(dbg_0.UNUSED_eu_mab_9_ ),
    .Y(_04214_)
  );
  INVX1 _11132_ (
    .A(dbg_0.UNUSED_eu_mab_8_ ),
    .Y(_04215_)
  );
  INVX1 _11133_ (
    .A(dbg_0.UNUSED_eu_mab_7_ ),
    .Y(_04216_)
  );
  INVX1 _11134_ (
    .A(dbg_0.UNUSED_eu_mab_6_ ),
    .Y(_04217_)
  );
  INVX1 _11135_ (
    .A(dbg_0.UNUSED_eu_mab_5_ ),
    .Y(_04218_)
  );
  INVX1 _11136_ (
    .A(dbg_0.UNUSED_eu_mab_4_ ),
    .Y(_04219_)
  );
  INVX1 _11137_ (
    .A(dbg_0.UNUSED_eu_mab_3_ ),
    .Y(_04220_)
  );
  INVX1 _11138_ (
    .A(dbg_0.UNUSED_eu_mab_2_ ),
    .Y(_04221_)
  );
  INVX1 _11139_ (
    .A(dbg_0.UNUSED_eu_mab_1_ ),
    .Y(_04222_)
  );
  INVX1 _11140_ (
    .A(_00144_),
    .Y(_04223_)
  );
  INVX1 _11141_ (
    .A(eu_mdb_out_0_),
    .Y(_04224_)
  );
  INVX1 _11142_ (
    .A(_00151_),
    .Y(_04225_)
  );
  INVX1 _11143_ (
    .A(eu_mdb_out_1_),
    .Y(_04226_)
  );
  INVX1 _11144_ (
    .A(_00152_),
    .Y(_04227_)
  );
  INVX1 _11145_ (
    .A(eu_mdb_out_2_),
    .Y(_04228_)
  );
  INVX1 _11146_ (
    .A(_00153_),
    .Y(_04229_)
  );
  INVX1 _11147_ (
    .A(eu_mdb_out_3_),
    .Y(_04230_)
  );
  INVX1 _11148_ (
    .A(_00154_),
    .Y(_04231_)
  );
  INVX1 _11149_ (
    .A(eu_mdb_out_4_),
    .Y(_04232_)
  );
  INVX1 _11150_ (
    .A(_00155_),
    .Y(_04233_)
  );
  INVX1 _11151_ (
    .A(eu_mdb_out_5_),
    .Y(_04234_)
  );
  INVX1 _11152_ (
    .A(_00156_),
    .Y(_04235_)
  );
  INVX1 _11153_ (
    .A(eu_mdb_out_6_),
    .Y(_04236_)
  );
  INVX1 _11154_ (
    .A(_00157_),
    .Y(_04237_)
  );
  INVX1 _11155_ (
    .A(eu_mdb_out_7_),
    .Y(_04238_)
  );
  INVX1 _11156_ (
    .A(_00158_),
    .Y(_04239_)
  );
  INVX1 _11157_ (
    .A(eu_mdb_out_8_),
    .Y(_04240_)
  );
  INVX1 _11158_ (
    .A(_00159_),
    .Y(_04241_)
  );
  INVX1 _11159_ (
    .A(eu_mdb_out_9_),
    .Y(_04242_)
  );
  INVX1 _11160_ (
    .A(_00145_),
    .Y(_04243_)
  );
  INVX1 _11161_ (
    .A(eu_mdb_out_10_),
    .Y(_04244_)
  );
  INVX1 _11162_ (
    .A(_00146_),
    .Y(_04245_)
  );
  INVX1 _11163_ (
    .A(eu_mdb_out_11_),
    .Y(_04246_)
  );
  INVX1 _11164_ (
    .A(_00147_),
    .Y(_04247_)
  );
  INVX1 _11165_ (
    .A(eu_mdb_out_12_),
    .Y(_04248_)
  );
  INVX1 _11166_ (
    .A(_00148_),
    .Y(_04249_)
  );
  INVX1 _11167_ (
    .A(eu_mdb_out_13_),
    .Y(_04250_)
  );
  INVX1 _11168_ (
    .A(_00149_),
    .Y(_04251_)
  );
  INVX1 _11169_ (
    .A(eu_mdb_out_14_),
    .Y(_04252_)
  );
  INVX1 _11170_ (
    .A(_00150_),
    .Y(_04253_)
  );
  INVX1 _11171_ (
    .A(eu_mdb_out_15_),
    .Y(_04254_)
  );
  INVX1 _11172_ (
    .A(dbg_0.UNUSED_eu_mb_wr_0_ ),
    .Y(_04255_)
  );
  INVX1 _11173_ (
    .A(dbg_0.dbg_mem_wr_0_ ),
    .Y(_04256_)
  );
  INVX1 _11174_ (
    .A(pmem_dout_0_),
    .Y(_04257_)
  );
  INVX1 _11175_ (
    .A(pmem_dout_1_),
    .Y(_04258_)
  );
  INVX1 _11176_ (
    .A(pmem_dout_2_),
    .Y(_04259_)
  );
  INVX1 _11177_ (
    .A(pmem_dout_3_),
    .Y(_04260_)
  );
  INVX1 _11178_ (
    .A(pmem_dout_4_),
    .Y(_04261_)
  );
  INVX1 _11179_ (
    .A(pmem_dout_5_),
    .Y(_04262_)
  );
  INVX1 _11180_ (
    .A(pmem_dout_6_),
    .Y(_04263_)
  );
  INVX1 _11181_ (
    .A(pmem_dout_7_),
    .Y(_04264_)
  );
  INVX1 _11182_ (
    .A(pmem_dout_8_),
    .Y(_04265_)
  );
  INVX1 _11183_ (
    .A(pmem_dout_9_),
    .Y(_04266_)
  );
  INVX1 _11184_ (
    .A(pmem_dout_10_),
    .Y(_04267_)
  );
  INVX1 _11185_ (
    .A(pmem_dout_11_),
    .Y(_04268_)
  );
  INVX1 _11186_ (
    .A(pmem_dout_12_),
    .Y(_04269_)
  );
  INVX1 _11187_ (
    .A(pmem_dout_13_),
    .Y(_04270_)
  );
  INVX1 _11188_ (
    .A(pmem_dout_14_),
    .Y(_04271_)
  );
  INVX1 _11189_ (
    .A(pmem_dout_15_),
    .Y(_04272_)
  );
  INVX1 _11190_ (
    .A(cpu_halt_st),
    .Y(_04273_)
  );
  INVX1 _11191_ (
    .A(_00162_),
    .Y(_04191_)
  );
  NOR2X1 _11192_ (
    .A(_04209_),
    .B(dbg_0.UNUSED_eu_mab_15_ ),
    .Y(_04274_)
  );
  INVX1 _11193_ (
    .A(_04274_),
    .Y(_04275_)
  );
  NAND3X1 _11194_ (
    .A(_04194_),
    .B(dbg_0.dbg_mem_addr_14_ ),
    .C(dbg_0.dbg_mem_en ),
    .Y(_04276_)
  );
  INVX1 _11195_ (
    .A(_04276_),
    .Y(_04277_)
  );
  AOI21X1 _11196_ (
    .A(dbg_0.UNUSED_eu_mab_14_ ),
    .B(_04274_),
    .C(_04276_),
    .Y(_04278_)
  );
  MUX2X1 _11197_ (
    .A(dbg_0.dbg_mem_wr_1_ ),
    .B(dbg_0.UNUSED_eu_mb_wr_1_ ),
    .S(_04278_),
    .Y(_00082_)
  );
  MUX2X1 _11198_ (
    .A(_04208_),
    .B(_04222_),
    .S(_04278_),
    .Y(_00051_)
  );
  MUX2X1 _11199_ (
    .A(_04207_),
    .B(_04221_),
    .S(_04278_),
    .Y(_00055_)
  );
  MUX2X1 _11200_ (
    .A(_04206_),
    .B(_04220_),
    .S(_04278_),
    .Y(_00056_)
  );
  MUX2X1 _11201_ (
    .A(_04205_),
    .B(_04219_),
    .S(_04278_),
    .Y(_00057_)
  );
  MUX2X1 _11202_ (
    .A(_04204_),
    .B(_04218_),
    .S(_04278_),
    .Y(_00058_)
  );
  MUX2X1 _11203_ (
    .A(_04203_),
    .B(_04217_),
    .S(_04278_),
    .Y(_00059_)
  );
  MUX2X1 _11204_ (
    .A(_04202_),
    .B(_04216_),
    .S(_04278_),
    .Y(_00060_)
  );
  MUX2X1 _11205_ (
    .A(_04201_),
    .B(_04215_),
    .S(_04278_),
    .Y(_00061_)
  );
  MUX2X1 _11206_ (
    .A(_04200_),
    .B(_04214_),
    .S(_04278_),
    .Y(_00062_)
  );
  MUX2X1 _11207_ (
    .A(_04199_),
    .B(_04213_),
    .S(_04278_),
    .Y(_00063_)
  );
  MUX2X1 _11208_ (
    .A(_04198_),
    .B(_04212_),
    .S(_04278_),
    .Y(_00052_)
  );
  MUX2X1 _11209_ (
    .A(_04197_),
    .B(_04211_),
    .S(_04278_),
    .Y(_00053_)
  );
  MUX2X1 _11210_ (
    .A(_04196_),
    .B(_04210_),
    .S(_04278_),
    .Y(_00054_)
  );
  MUX2X1 _11211_ (
    .A(_04223_),
    .B(_04224_),
    .S(_04278_),
    .Y(_00065_)
  );
  MUX2X1 _11212_ (
    .A(_04225_),
    .B(_04226_),
    .S(_04278_),
    .Y(_00072_)
  );
  MUX2X1 _11213_ (
    .A(_04227_),
    .B(_04228_),
    .S(_04278_),
    .Y(_00073_)
  );
  MUX2X1 _11214_ (
    .A(_04229_),
    .B(_04230_),
    .S(_04278_),
    .Y(_00074_)
  );
  MUX2X1 _11215_ (
    .A(_04231_),
    .B(_04232_),
    .S(_04278_),
    .Y(_00075_)
  );
  MUX2X1 _11216_ (
    .A(_04233_),
    .B(_04234_),
    .S(_04278_),
    .Y(_00076_)
  );
  MUX2X1 _11217_ (
    .A(_04235_),
    .B(_04236_),
    .S(_04278_),
    .Y(_00077_)
  );
  MUX2X1 _11218_ (
    .A(_04237_),
    .B(_04238_),
    .S(_04278_),
    .Y(_00078_)
  );
  MUX2X1 _11219_ (
    .A(_04239_),
    .B(_04240_),
    .S(_04278_),
    .Y(_00079_)
  );
  MUX2X1 _11220_ (
    .A(_04241_),
    .B(_04242_),
    .S(_04278_),
    .Y(_00080_)
  );
  MUX2X1 _11221_ (
    .A(_04243_),
    .B(_04244_),
    .S(_04278_),
    .Y(_00066_)
  );
  MUX2X1 _11222_ (
    .A(_04245_),
    .B(_04246_),
    .S(_04278_),
    .Y(_00067_)
  );
  MUX2X1 _11223_ (
    .A(_04247_),
    .B(_04248_),
    .S(_04278_),
    .Y(_00068_)
  );
  MUX2X1 _11224_ (
    .A(_04249_),
    .B(_04250_),
    .S(_04278_),
    .Y(_00069_)
  );
  MUX2X1 _11225_ (
    .A(_04251_),
    .B(_04252_),
    .S(_04278_),
    .Y(_00070_)
  );
  MUX2X1 _11226_ (
    .A(_04253_),
    .B(_04254_),
    .S(_04278_),
    .Y(_00071_)
  );
  OR2X1 _11227_ (
    .A(dbg_0.UNUSED_eu_mb_wr_1_ ),
    .B(dbg_0.UNUSED_eu_mb_wr_0_ ),
    .Y(_04279_)
  );
  NAND2X1 _11228_ (
    .A(dbg_0.UNUSED_eu_mb_en ),
    .B(dbg_0.UNUSED_eu_mab_15_ ),
    .Y(_04280_)
  );
  NOR2X1 _11229_ (
    .A(_04279_),
    .B(_04280_),
    .Y(mem_backbone_0.eu_pmem_en )
  );
  NAND2X1 _11230_ (
    .A(execution_unit_0.pc_nxt_15_ ),
    .B(fe_mb_en),
    .Y(_04281_)
  );
  INVX1 _11231_ (
    .A(_04281_),
    .Y(mem_backbone_0.fe_pmem_en )
  );
  OAI21X1 _11232_ (
    .A(_04279_),
    .B(_04280_),
    .C(_04281_),
    .Y(_04282_)
  );
  NAND2X1 _11233_ (
    .A(dbg_0.dbg_mem_addr_15_ ),
    .B(dbg_0.dbg_mem_en ),
    .Y(_04283_)
  );
  NOR2X1 _11234_ (
    .A(_04282_),
    .B(_04283_),
    .Y(mem_backbone_0.ext_pmem_en )
  );
  NAND2X1 _11235_ (
    .A(dbg_0.dbg_mem_wr_0_ ),
    .B(mem_backbone_0.ext_pmem_en ),
    .Y(_00160_)
  );
  NAND2X1 _11236_ (
    .A(dbg_0.dbg_mem_wr_1_ ),
    .B(mem_backbone_0.ext_pmem_en ),
    .Y(_00161_)
  );
  MUX2X1 _11237_ (
    .A(dbg_0.UNUSED_eu_mab_1_ ),
    .B(execution_unit_0.pc_nxt_1_ ),
    .S(mem_backbone_0.eu_pmem_en ),
    .Y(_04284_)
  );
  MUX2X1 _11238_ (
    .A(_04208_),
    .B(_04284_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00129_)
  );
  MUX2X1 _11239_ (
    .A(dbg_0.UNUSED_eu_mab_2_ ),
    .B(execution_unit_0.pc_nxt_2_ ),
    .S(mem_backbone_0.eu_pmem_en ),
    .Y(_04285_)
  );
  MUX2X1 _11240_ (
    .A(_04207_),
    .B(_04285_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00134_)
  );
  MUX2X1 _11241_ (
    .A(dbg_0.UNUSED_eu_mab_3_ ),
    .B(execution_unit_0.pc_nxt_3_ ),
    .S(mem_backbone_0.eu_pmem_en ),
    .Y(_04286_)
  );
  MUX2X1 _11242_ (
    .A(_04206_),
    .B(_04286_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00135_)
  );
  MUX2X1 _11243_ (
    .A(dbg_0.UNUSED_eu_mab_4_ ),
    .B(execution_unit_0.pc_nxt_4_ ),
    .S(mem_backbone_0.eu_pmem_en ),
    .Y(_04287_)
  );
  MUX2X1 _11244_ (
    .A(_04205_),
    .B(_04287_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00136_)
  );
  MUX2X1 _11245_ (
    .A(dbg_0.UNUSED_eu_mab_5_ ),
    .B(execution_unit_0.pc_nxt_5_ ),
    .S(mem_backbone_0.eu_pmem_en ),
    .Y(_04288_)
  );
  MUX2X1 _11246_ (
    .A(_04204_),
    .B(_04288_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00137_)
  );
  MUX2X1 _11247_ (
    .A(dbg_0.UNUSED_eu_mab_6_ ),
    .B(execution_unit_0.pc_nxt_6_ ),
    .S(mem_backbone_0.eu_pmem_en ),
    .Y(_04289_)
  );
  MUX2X1 _11248_ (
    .A(_04203_),
    .B(_04289_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00138_)
  );
  MUX2X1 _11249_ (
    .A(dbg_0.UNUSED_eu_mab_7_ ),
    .B(execution_unit_0.pc_nxt_7_ ),
    .S(mem_backbone_0.eu_pmem_en ),
    .Y(_04290_)
  );
  MUX2X1 _11250_ (
    .A(_04202_),
    .B(_04290_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00139_)
  );
  MUX2X1 _11251_ (
    .A(dbg_0.UNUSED_eu_mab_8_ ),
    .B(execution_unit_0.pc_nxt_8_ ),
    .S(mem_backbone_0.eu_pmem_en ),
    .Y(_04291_)
  );
  MUX2X1 _11252_ (
    .A(_04201_),
    .B(_04291_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00140_)
  );
  MUX2X1 _11253_ (
    .A(dbg_0.UNUSED_eu_mab_9_ ),
    .B(execution_unit_0.pc_nxt_9_ ),
    .S(mem_backbone_0.eu_pmem_en ),
    .Y(_04292_)
  );
  MUX2X1 _11254_ (
    .A(_04200_),
    .B(_04292_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00141_)
  );
  MUX2X1 _11255_ (
    .A(dbg_0.UNUSED_eu_mab_10_ ),
    .B(execution_unit_0.pc_nxt_10_ ),
    .S(mem_backbone_0.eu_pmem_en ),
    .Y(_04293_)
  );
  MUX2X1 _11256_ (
    .A(_04199_),
    .B(_04293_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00142_)
  );
  MUX2X1 _11257_ (
    .A(dbg_0.UNUSED_eu_mab_11_ ),
    .B(execution_unit_0.pc_nxt_11_ ),
    .S(mem_backbone_0.eu_pmem_en ),
    .Y(_04294_)
  );
  MUX2X1 _11258_ (
    .A(_04198_),
    .B(_04294_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00130_)
  );
  MUX2X1 _11259_ (
    .A(dbg_0.UNUSED_eu_mab_12_ ),
    .B(execution_unit_0.pc_nxt_12_ ),
    .S(mem_backbone_0.eu_pmem_en ),
    .Y(_04295_)
  );
  MUX2X1 _11260_ (
    .A(_04197_),
    .B(_04295_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00131_)
  );
  MUX2X1 _11261_ (
    .A(dbg_0.UNUSED_eu_mab_13_ ),
    .B(execution_unit_0.pc_nxt_13_ ),
    .S(mem_backbone_0.eu_pmem_en ),
    .Y(_04296_)
  );
  MUX2X1 _11262_ (
    .A(_04196_),
    .B(_04296_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00132_)
  );
  MUX2X1 _11263_ (
    .A(dbg_0.UNUSED_eu_mab_14_ ),
    .B(execution_unit_0.pc_nxt_14_ ),
    .S(mem_backbone_0.eu_pmem_en ),
    .Y(_04297_)
  );
  MUX2X1 _11264_ (
    .A(_04195_),
    .B(_04297_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00133_)
  );
  NOR3X1 _11265_ (
    .A(_04209_),
    .B(dbg_0.UNUSED_eu_mab_15_ ),
    .C(dbg_0.UNUSED_eu_mab_14_ ),
    .Y(mem_backbone_0.eu_per_en )
  );
  NAND3X1 _11266_ (
    .A(_04194_),
    .B(_04195_),
    .C(dbg_0.dbg_mem_en ),
    .Y(_04298_)
  );
  NOR2X1 _11267_ (
    .A(mem_backbone_0.eu_per_en ),
    .B(_04298_),
    .Y(mem_backbone_0.ext_per_en )
  );
  MUX2X1 _11268_ (
    .A(_04256_),
    .B(_04255_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00127_)
  );
  MUX2X1 _11269_ (
    .A(_04193_),
    .B(_04192_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00128_)
  );
  MUX2X1 _11270_ (
    .A(_04208_),
    .B(_04222_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00097_)
  );
  MUX2X1 _11271_ (
    .A(_04207_),
    .B(_04221_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00101_)
  );
  MUX2X1 _11272_ (
    .A(_04206_),
    .B(_04220_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00102_)
  );
  MUX2X1 _11273_ (
    .A(_04205_),
    .B(_04219_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00103_)
  );
  MUX2X1 _11274_ (
    .A(_04204_),
    .B(_04218_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00104_)
  );
  MUX2X1 _11275_ (
    .A(_04203_),
    .B(_04217_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00105_)
  );
  MUX2X1 _11276_ (
    .A(_04202_),
    .B(_04216_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00106_)
  );
  MUX2X1 _11277_ (
    .A(_04201_),
    .B(_04215_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00107_)
  );
  MUX2X1 _11278_ (
    .A(_04200_),
    .B(_04214_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00108_)
  );
  MUX2X1 _11279_ (
    .A(_04199_),
    .B(_04213_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00109_)
  );
  MUX2X1 _11280_ (
    .A(_04198_),
    .B(_04212_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00098_)
  );
  MUX2X1 _11281_ (
    .A(_04197_),
    .B(_04211_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00099_)
  );
  MUX2X1 _11282_ (
    .A(_04196_),
    .B(_04210_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00100_)
  );
  MUX2X1 _11283_ (
    .A(_04223_),
    .B(_04224_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00110_)
  );
  MUX2X1 _11284_ (
    .A(_04225_),
    .B(_04226_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00117_)
  );
  MUX2X1 _11285_ (
    .A(_04227_),
    .B(_04228_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00118_)
  );
  MUX2X1 _11286_ (
    .A(_04229_),
    .B(_04230_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00119_)
  );
  MUX2X1 _11287_ (
    .A(_04231_),
    .B(_04232_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00120_)
  );
  MUX2X1 _11288_ (
    .A(_04233_),
    .B(_04234_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00121_)
  );
  MUX2X1 _11289_ (
    .A(_04235_),
    .B(_04236_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00122_)
  );
  MUX2X1 _11290_ (
    .A(_04237_),
    .B(_04238_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00123_)
  );
  MUX2X1 _11291_ (
    .A(_04239_),
    .B(_04240_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00124_)
  );
  MUX2X1 _11292_ (
    .A(_04241_),
    .B(_04242_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00125_)
  );
  MUX2X1 _11293_ (
    .A(_04243_),
    .B(_04244_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00111_)
  );
  MUX2X1 _11294_ (
    .A(_04245_),
    .B(_04246_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00112_)
  );
  MUX2X1 _11295_ (
    .A(_04247_),
    .B(_04248_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00113_)
  );
  MUX2X1 _11296_ (
    .A(_04249_),
    .B(_04250_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00114_)
  );
  MUX2X1 _11297_ (
    .A(_04251_),
    .B(_04252_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00115_)
  );
  MUX2X1 _11298_ (
    .A(_04253_),
    .B(_04254_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00116_)
  );
  NAND2X1 _11299_ (
    .A(mem_backbone_0.pmem_dout_bckup_0_ ),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04299_)
  );
  OAI21X1 _11300_ (
    .A(_04257_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04299_),
    .Y(dbg_0.fe_mdb_in_0_ )
  );
  NAND2X1 _11301_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_1_ ),
    .Y(_04300_)
  );
  OAI21X1 _11302_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04258_),
    .C(_04300_),
    .Y(dbg_0.fe_mdb_in_1_ )
  );
  NAND2X1 _11303_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_2_ ),
    .Y(_04301_)
  );
  OAI21X1 _11304_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04259_),
    .C(_04301_),
    .Y(dbg_0.fe_mdb_in_2_ )
  );
  NAND2X1 _11305_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_3_ ),
    .Y(_04302_)
  );
  OAI21X1 _11306_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04260_),
    .C(_04302_),
    .Y(dbg_0.fe_mdb_in_3_ )
  );
  NAND2X1 _11307_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_4_ ),
    .Y(_04303_)
  );
  OAI21X1 _11308_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04261_),
    .C(_04303_),
    .Y(dbg_0.fe_mdb_in_4_ )
  );
  NAND2X1 _11309_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_5_ ),
    .Y(_04304_)
  );
  OAI21X1 _11310_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04262_),
    .C(_04304_),
    .Y(dbg_0.fe_mdb_in_5_ )
  );
  NAND2X1 _11311_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_6_ ),
    .Y(_04305_)
  );
  OAI21X1 _11312_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04263_),
    .C(_04305_),
    .Y(dbg_0.fe_mdb_in_6_ )
  );
  NAND2X1 _11313_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_7_ ),
    .Y(_04306_)
  );
  OAI21X1 _11314_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04264_),
    .C(_04306_),
    .Y(dbg_0.fe_mdb_in_7_ )
  );
  NAND2X1 _11315_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_8_ ),
    .Y(_04307_)
  );
  OAI21X1 _11316_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04265_),
    .C(_04307_),
    .Y(dbg_0.fe_mdb_in_8_ )
  );
  NAND2X1 _11317_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_9_ ),
    .Y(_04308_)
  );
  OAI21X1 _11318_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04266_),
    .C(_04308_),
    .Y(dbg_0.fe_mdb_in_9_ )
  );
  NAND2X1 _11319_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_10_ ),
    .Y(_04309_)
  );
  OAI21X1 _11320_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04267_),
    .C(_04309_),
    .Y(dbg_0.fe_mdb_in_10_ )
  );
  NAND2X1 _11321_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_11_ ),
    .Y(_04310_)
  );
  OAI21X1 _11322_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04268_),
    .C(_04310_),
    .Y(dbg_0.fe_mdb_in_11_ )
  );
  NAND2X1 _11323_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_12_ ),
    .Y(_04311_)
  );
  OAI21X1 _11324_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04269_),
    .C(_04311_),
    .Y(dbg_0.fe_mdb_in_12_ )
  );
  NAND2X1 _11325_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_13_ ),
    .Y(_04312_)
  );
  OAI21X1 _11326_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04270_),
    .C(_04312_),
    .Y(dbg_0.fe_mdb_in_13_ )
  );
  NAND2X1 _11327_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_14_ ),
    .Y(_04313_)
  );
  OAI21X1 _11328_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04271_),
    .C(_04313_),
    .Y(dbg_0.fe_mdb_in_14_ )
  );
  NAND2X1 _11329_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(mem_backbone_0.pmem_dout_bckup_15_ ),
    .Y(_04314_)
  );
  OAI21X1 _11330_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04272_),
    .C(_04314_),
    .Y(dbg_0.fe_mdb_in_15_ )
  );
  MUX2X1 _11331_ (
    .A(mem_backbone_0.per_dout_val_0_ ),
    .B(dmem_dout_0_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04315_)
  );
  NAND2X1 _11332_ (
    .A(pmem_dout_0_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04316_)
  );
  OAI21X1 _11333_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04315_),
    .C(_04316_),
    .Y(eu_mdb_in_0_)
  );
  MUX2X1 _11334_ (
    .A(mem_backbone_0.per_dout_val_1_ ),
    .B(dmem_dout_1_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04317_)
  );
  NAND2X1 _11335_ (
    .A(pmem_dout_1_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04318_)
  );
  OAI21X1 _11336_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04317_),
    .C(_04318_),
    .Y(eu_mdb_in_1_)
  );
  MUX2X1 _11337_ (
    .A(mem_backbone_0.per_dout_val_2_ ),
    .B(dmem_dout_2_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04319_)
  );
  NAND2X1 _11338_ (
    .A(pmem_dout_2_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04320_)
  );
  OAI21X1 _11339_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04319_),
    .C(_04320_),
    .Y(eu_mdb_in_2_)
  );
  MUX2X1 _11340_ (
    .A(mem_backbone_0.per_dout_val_3_ ),
    .B(dmem_dout_3_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04321_)
  );
  NAND2X1 _11341_ (
    .A(pmem_dout_3_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04322_)
  );
  OAI21X1 _11342_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04321_),
    .C(_04322_),
    .Y(eu_mdb_in_3_)
  );
  MUX2X1 _11343_ (
    .A(mem_backbone_0.per_dout_val_4_ ),
    .B(dmem_dout_4_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04323_)
  );
  NAND2X1 _11344_ (
    .A(pmem_dout_4_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04324_)
  );
  OAI21X1 _11345_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04323_),
    .C(_04324_),
    .Y(eu_mdb_in_4_)
  );
  MUX2X1 _11346_ (
    .A(mem_backbone_0.per_dout_val_5_ ),
    .B(dmem_dout_5_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04325_)
  );
  NAND2X1 _11347_ (
    .A(pmem_dout_5_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04326_)
  );
  OAI21X1 _11348_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04325_),
    .C(_04326_),
    .Y(eu_mdb_in_5_)
  );
  MUX2X1 _11349_ (
    .A(mem_backbone_0.per_dout_val_6_ ),
    .B(dmem_dout_6_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04327_)
  );
  NAND2X1 _11350_ (
    .A(pmem_dout_6_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04328_)
  );
  OAI21X1 _11351_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04327_),
    .C(_04328_),
    .Y(eu_mdb_in_6_)
  );
  MUX2X1 _11352_ (
    .A(mem_backbone_0.per_dout_val_7_ ),
    .B(dmem_dout_7_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04329_)
  );
  NAND2X1 _11353_ (
    .A(pmem_dout_7_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04330_)
  );
  OAI21X1 _11354_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04329_),
    .C(_04330_),
    .Y(eu_mdb_in_7_)
  );
  MUX2X1 _11355_ (
    .A(mem_backbone_0.per_dout_val_8_ ),
    .B(dmem_dout_8_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04331_)
  );
  NAND2X1 _11356_ (
    .A(pmem_dout_8_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04332_)
  );
  OAI21X1 _11357_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04331_),
    .C(_04332_),
    .Y(eu_mdb_in_8_)
  );
  MUX2X1 _11358_ (
    .A(mem_backbone_0.per_dout_val_9_ ),
    .B(dmem_dout_9_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04333_)
  );
  NAND2X1 _11359_ (
    .A(pmem_dout_9_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04334_)
  );
  OAI21X1 _11360_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04333_),
    .C(_04334_),
    .Y(eu_mdb_in_9_)
  );
  MUX2X1 _11361_ (
    .A(mem_backbone_0.per_dout_val_10_ ),
    .B(dmem_dout_10_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04335_)
  );
  NAND2X1 _11362_ (
    .A(pmem_dout_10_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04336_)
  );
  OAI21X1 _11363_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04335_),
    .C(_04336_),
    .Y(eu_mdb_in_10_)
  );
  MUX2X1 _11364_ (
    .A(mem_backbone_0.per_dout_val_11_ ),
    .B(dmem_dout_11_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04337_)
  );
  NAND2X1 _11365_ (
    .A(pmem_dout_11_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04338_)
  );
  OAI21X1 _11366_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04337_),
    .C(_04338_),
    .Y(eu_mdb_in_11_)
  );
  MUX2X1 _11367_ (
    .A(mem_backbone_0.per_dout_val_12_ ),
    .B(dmem_dout_12_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04339_)
  );
  NAND2X1 _11368_ (
    .A(pmem_dout_12_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04340_)
  );
  OAI21X1 _11369_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04339_),
    .C(_04340_),
    .Y(eu_mdb_in_12_)
  );
  MUX2X1 _11370_ (
    .A(mem_backbone_0.per_dout_val_13_ ),
    .B(dmem_dout_13_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04341_)
  );
  NAND2X1 _11371_ (
    .A(pmem_dout_13_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04342_)
  );
  OAI21X1 _11372_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04341_),
    .C(_04342_),
    .Y(eu_mdb_in_13_)
  );
  MUX2X1 _11373_ (
    .A(mem_backbone_0.per_dout_val_14_ ),
    .B(dmem_dout_14_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04343_)
  );
  NAND2X1 _11374_ (
    .A(pmem_dout_14_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04344_)
  );
  OAI21X1 _11375_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04343_),
    .C(_04344_),
    .Y(eu_mdb_in_14_)
  );
  MUX2X1 _11376_ (
    .A(mem_backbone_0.per_dout_val_15_ ),
    .B(dmem_dout_15_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04345_)
  );
  NAND2X1 _11377_ (
    .A(pmem_dout_15_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04346_)
  );
  OAI21X1 _11378_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04345_),
    .C(_04346_),
    .Y(eu_mdb_in_15_)
  );
  MUX2X1 _11379_ (
    .A(mem_backbone_0.per_dout_val_0_ ),
    .B(dmem_dout_0_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04347_)
  );
  NAND2X1 _11380_ (
    .A(pmem_dout_0_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04348_)
  );
  OAI21X1 _11381_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04347_),
    .C(_04348_),
    .Y(dbg_0.dbg_mem_din_0_ )
  );
  MUX2X1 _11382_ (
    .A(mem_backbone_0.per_dout_val_1_ ),
    .B(dmem_dout_1_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04349_)
  );
  NAND2X1 _11383_ (
    .A(pmem_dout_1_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04350_)
  );
  OAI21X1 _11384_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04349_),
    .C(_04350_),
    .Y(dbg_0.dbg_mem_din_1_ )
  );
  MUX2X1 _11385_ (
    .A(mem_backbone_0.per_dout_val_2_ ),
    .B(dmem_dout_2_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04351_)
  );
  NAND2X1 _11386_ (
    .A(pmem_dout_2_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04352_)
  );
  OAI21X1 _11387_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04351_),
    .C(_04352_),
    .Y(dbg_0.dbg_mem_din_2_ )
  );
  MUX2X1 _11388_ (
    .A(mem_backbone_0.per_dout_val_3_ ),
    .B(dmem_dout_3_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04353_)
  );
  NAND2X1 _11389_ (
    .A(pmem_dout_3_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04354_)
  );
  OAI21X1 _11390_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04353_),
    .C(_04354_),
    .Y(dbg_0.dbg_mem_din_3_ )
  );
  MUX2X1 _11391_ (
    .A(mem_backbone_0.per_dout_val_4_ ),
    .B(dmem_dout_4_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04355_)
  );
  NAND2X1 _11392_ (
    .A(pmem_dout_4_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04356_)
  );
  OAI21X1 _11393_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04355_),
    .C(_04356_),
    .Y(dbg_0.dbg_mem_din_4_ )
  );
  MUX2X1 _11394_ (
    .A(mem_backbone_0.per_dout_val_5_ ),
    .B(dmem_dout_5_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04357_)
  );
  NAND2X1 _11395_ (
    .A(pmem_dout_5_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04358_)
  );
  OAI21X1 _11396_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04357_),
    .C(_04358_),
    .Y(dbg_0.dbg_mem_din_5_ )
  );
  MUX2X1 _11397_ (
    .A(mem_backbone_0.per_dout_val_6_ ),
    .B(dmem_dout_6_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04359_)
  );
  NAND2X1 _11398_ (
    .A(pmem_dout_6_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04360_)
  );
  OAI21X1 _11399_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04359_),
    .C(_04360_),
    .Y(dbg_0.dbg_mem_din_6_ )
  );
  MUX2X1 _11400_ (
    .A(mem_backbone_0.per_dout_val_7_ ),
    .B(dmem_dout_7_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04361_)
  );
  NAND2X1 _11401_ (
    .A(pmem_dout_7_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04362_)
  );
  OAI21X1 _11402_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04361_),
    .C(_04362_),
    .Y(dbg_0.dbg_mem_din_7_ )
  );
  MUX2X1 _11403_ (
    .A(mem_backbone_0.per_dout_val_8_ ),
    .B(dmem_dout_8_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04363_)
  );
  NAND2X1 _11404_ (
    .A(pmem_dout_8_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04364_)
  );
  OAI21X1 _11405_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04363_),
    .C(_04364_),
    .Y(dbg_0.dbg_mem_din_8_ )
  );
  MUX2X1 _11406_ (
    .A(mem_backbone_0.per_dout_val_9_ ),
    .B(dmem_dout_9_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04365_)
  );
  NAND2X1 _11407_ (
    .A(pmem_dout_9_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04366_)
  );
  OAI21X1 _11408_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04365_),
    .C(_04366_),
    .Y(dbg_0.dbg_mem_din_9_ )
  );
  MUX2X1 _11409_ (
    .A(mem_backbone_0.per_dout_val_10_ ),
    .B(dmem_dout_10_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04367_)
  );
  NAND2X1 _11410_ (
    .A(pmem_dout_10_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04368_)
  );
  OAI21X1 _11411_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04367_),
    .C(_04368_),
    .Y(dbg_0.dbg_mem_din_10_ )
  );
  MUX2X1 _11412_ (
    .A(mem_backbone_0.per_dout_val_11_ ),
    .B(dmem_dout_11_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04369_)
  );
  NAND2X1 _11413_ (
    .A(pmem_dout_11_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04370_)
  );
  OAI21X1 _11414_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04369_),
    .C(_04370_),
    .Y(dbg_0.dbg_mem_din_11_ )
  );
  MUX2X1 _11415_ (
    .A(mem_backbone_0.per_dout_val_12_ ),
    .B(dmem_dout_12_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04371_)
  );
  NAND2X1 _11416_ (
    .A(pmem_dout_12_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04372_)
  );
  OAI21X1 _11417_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04371_),
    .C(_04372_),
    .Y(dbg_0.dbg_mem_din_12_ )
  );
  MUX2X1 _11418_ (
    .A(mem_backbone_0.per_dout_val_13_ ),
    .B(dmem_dout_13_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04373_)
  );
  NAND2X1 _11419_ (
    .A(pmem_dout_13_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04374_)
  );
  OAI21X1 _11420_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04373_),
    .C(_04374_),
    .Y(dbg_0.dbg_mem_din_13_ )
  );
  MUX2X1 _11421_ (
    .A(mem_backbone_0.per_dout_val_14_ ),
    .B(dmem_dout_14_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04375_)
  );
  NAND2X1 _11422_ (
    .A(pmem_dout_14_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04376_)
  );
  OAI21X1 _11423_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04375_),
    .C(_04376_),
    .Y(dbg_0.dbg_mem_din_14_ )
  );
  MUX2X1 _11424_ (
    .A(mem_backbone_0.per_dout_val_15_ ),
    .B(dmem_dout_15_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04377_)
  );
  NAND2X1 _11425_ (
    .A(pmem_dout_15_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04378_)
  );
  OAI21X1 _11426_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04377_),
    .C(_04378_),
    .Y(dbg_0.dbg_mem_din_15_ )
  );
  NAND3X1 _11427_ (
    .A(_04273_),
    .B(mem_backbone_0.fe_pmem_en_dly ),
    .C(_04281_),
    .Y(_04379_)
  );
  MUX2X1 _11428_ (
    .A(mem_backbone_0.pmem_dout_bckup_0_ ),
    .B(pmem_dout_0_),
    .S(_04379_),
    .Y(_04380_)
  );
  INVX1 _11429_ (
    .A(_04380_),
    .Y(_04174_)
  );
  MUX2X1 _11430_ (
    .A(mem_backbone_0.pmem_dout_bckup_1_ ),
    .B(pmem_dout_1_),
    .S(_04379_),
    .Y(_04381_)
  );
  INVX1 _11431_ (
    .A(_04381_),
    .Y(_04181_)
  );
  MUX2X1 _11432_ (
    .A(mem_backbone_0.pmem_dout_bckup_2_ ),
    .B(pmem_dout_2_),
    .S(_04379_),
    .Y(_04382_)
  );
  INVX1 _11433_ (
    .A(_04382_),
    .Y(_04182_)
  );
  MUX2X1 _11434_ (
    .A(mem_backbone_0.pmem_dout_bckup_3_ ),
    .B(pmem_dout_3_),
    .S(_04379_),
    .Y(_04383_)
  );
  INVX1 _11435_ (
    .A(_04383_),
    .Y(_04183_)
  );
  MUX2X1 _11436_ (
    .A(mem_backbone_0.pmem_dout_bckup_4_ ),
    .B(pmem_dout_4_),
    .S(_04379_),
    .Y(_04384_)
  );
  INVX1 _11437_ (
    .A(_04384_),
    .Y(_04184_)
  );
  MUX2X1 _11438_ (
    .A(mem_backbone_0.pmem_dout_bckup_5_ ),
    .B(pmem_dout_5_),
    .S(_04379_),
    .Y(_04385_)
  );
  INVX1 _11439_ (
    .A(_04385_),
    .Y(_04185_)
  );
  MUX2X1 _11440_ (
    .A(mem_backbone_0.pmem_dout_bckup_6_ ),
    .B(pmem_dout_6_),
    .S(_04379_),
    .Y(_04386_)
  );
  INVX1 _11441_ (
    .A(_04386_),
    .Y(_04186_)
  );
  MUX2X1 _11442_ (
    .A(mem_backbone_0.pmem_dout_bckup_7_ ),
    .B(pmem_dout_7_),
    .S(_04379_),
    .Y(_04387_)
  );
  INVX1 _11443_ (
    .A(_04387_),
    .Y(_04187_)
  );
  MUX2X1 _11444_ (
    .A(mem_backbone_0.pmem_dout_bckup_8_ ),
    .B(pmem_dout_8_),
    .S(_04379_),
    .Y(_04388_)
  );
  INVX1 _11445_ (
    .A(_04388_),
    .Y(_04188_)
  );
  MUX2X1 _11446_ (
    .A(mem_backbone_0.pmem_dout_bckup_9_ ),
    .B(pmem_dout_9_),
    .S(_04379_),
    .Y(_04389_)
  );
  INVX1 _11447_ (
    .A(_04389_),
    .Y(_04189_)
  );
  MUX2X1 _11448_ (
    .A(mem_backbone_0.pmem_dout_bckup_10_ ),
    .B(pmem_dout_10_),
    .S(_04379_),
    .Y(_04390_)
  );
  INVX1 _11449_ (
    .A(_04390_),
    .Y(_04175_)
  );
  MUX2X1 _11450_ (
    .A(mem_backbone_0.pmem_dout_bckup_11_ ),
    .B(pmem_dout_11_),
    .S(_04379_),
    .Y(_04391_)
  );
  INVX1 _11451_ (
    .A(_04391_),
    .Y(_04176_)
  );
  MUX2X1 _11452_ (
    .A(mem_backbone_0.pmem_dout_bckup_12_ ),
    .B(pmem_dout_12_),
    .S(_04379_),
    .Y(_04392_)
  );
  INVX1 _11453_ (
    .A(_04392_),
    .Y(_04177_)
  );
  MUX2X1 _11454_ (
    .A(mem_backbone_0.pmem_dout_bckup_13_ ),
    .B(pmem_dout_13_),
    .S(_04379_),
    .Y(_04393_)
  );
  INVX1 _11455_ (
    .A(_04393_),
    .Y(_04178_)
  );
  MUX2X1 _11456_ (
    .A(mem_backbone_0.pmem_dout_bckup_14_ ),
    .B(pmem_dout_14_),
    .S(_04379_),
    .Y(_04394_)
  );
  INVX1 _11457_ (
    .A(_04394_),
    .Y(_04179_)
  );
  MUX2X1 _11458_ (
    .A(mem_backbone_0.pmem_dout_bckup_15_ ),
    .B(pmem_dout_15_),
    .S(_04379_),
    .Y(_04395_)
  );
  INVX1 _11459_ (
    .A(_04395_),
    .Y(_04180_)
  );
  MUX2X1 _11460_ (
    .A(dbg_0.dbg_mem_wr_0_ ),
    .B(dbg_0.UNUSED_eu_mb_wr_0_ ),
    .S(_04278_),
    .Y(_00081_)
  );
  NOR2X1 _11461_ (
    .A(_04282_),
    .B(mem_backbone_0.ext_pmem_en ),
    .Y(_00143_)
  );
  AOI21X1 _11462_ (
    .A(dbg_0.UNUSED_eu_mab_14_ ),
    .B(_04274_),
    .C(_04277_),
    .Y(_00064_)
  );
  AND2X1 _11463_ (
    .A(mem_backbone_0.eu_pmem_en ),
    .B(mem_backbone_0.fe_pmem_en ),
    .Y(fe_pmem_wait)
  );
  OAI21X1 _11464_ (
    .A(dbg_0.UNUSED_eu_mab_14_ ),
    .B(_04275_),
    .C(_04298_),
    .Y(_00126_)
  );
  NOR2X1 _11465_ (
    .A(mem_backbone_0.fe_pmem_en_dly ),
    .B(_04281_),
    .Y(_04396_)
  );
  NAND2X1 _11466_ (
    .A(mem_backbone_0.pmem_dout_bckup_sel ),
    .B(_04273_),
    .Y(_04397_)
  );
  OAI21X1 _11467_ (
    .A(_04396_),
    .B(_04397_),
    .C(_04379_),
    .Y(_04190_)
  );
  DFFSR _11468_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.ext_per_en ),
    .Q(mem_backbone_0.ext_mem_din_sel_0_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11469_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.ext_pmem_en ),
    .Q(mem_backbone_0.ext_mem_din_sel_1_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11470_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.eu_per_en ),
    .Q(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11471_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.eu_pmem_en ),
    .Q(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11472_ (
    .CLK(dco_clk),
    .D(_04190_),
    .Q(mem_backbone_0.pmem_dout_bckup_sel ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11473_ (
    .CLK(dco_clk),
    .D(_04174_),
    .Q(mem_backbone_0.pmem_dout_bckup_0_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11474_ (
    .CLK(dco_clk),
    .D(_04181_),
    .Q(mem_backbone_0.pmem_dout_bckup_1_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11475_ (
    .CLK(dco_clk),
    .D(_04182_),
    .Q(mem_backbone_0.pmem_dout_bckup_2_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11476_ (
    .CLK(dco_clk),
    .D(_04183_),
    .Q(mem_backbone_0.pmem_dout_bckup_3_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11477_ (
    .CLK(dco_clk),
    .D(_04184_),
    .Q(mem_backbone_0.pmem_dout_bckup_4_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11478_ (
    .CLK(dco_clk),
    .D(_04185_),
    .Q(mem_backbone_0.pmem_dout_bckup_5_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11479_ (
    .CLK(dco_clk),
    .D(_04186_),
    .Q(mem_backbone_0.pmem_dout_bckup_6_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11480_ (
    .CLK(dco_clk),
    .D(_04187_),
    .Q(mem_backbone_0.pmem_dout_bckup_7_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11481_ (
    .CLK(dco_clk),
    .D(_04188_),
    .Q(mem_backbone_0.pmem_dout_bckup_8_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11482_ (
    .CLK(dco_clk),
    .D(_04189_),
    .Q(mem_backbone_0.pmem_dout_bckup_9_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11483_ (
    .CLK(dco_clk),
    .D(_04175_),
    .Q(mem_backbone_0.pmem_dout_bckup_10_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11484_ (
    .CLK(dco_clk),
    .D(_04176_),
    .Q(mem_backbone_0.pmem_dout_bckup_11_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11485_ (
    .CLK(dco_clk),
    .D(_04177_),
    .Q(mem_backbone_0.pmem_dout_bckup_12_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11486_ (
    .CLK(dco_clk),
    .D(_04178_),
    .Q(mem_backbone_0.pmem_dout_bckup_13_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11487_ (
    .CLK(dco_clk),
    .D(_04179_),
    .Q(mem_backbone_0.pmem_dout_bckup_14_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11488_ (
    .CLK(dco_clk),
    .D(_04180_),
    .Q(mem_backbone_0.pmem_dout_bckup_15_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11489_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.fe_pmem_en ),
    .Q(mem_backbone_0.fe_pmem_en_dly ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11490_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_0_ ),
    .Q(mem_backbone_0.per_dout_val_0_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11491_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_1_ ),
    .Q(mem_backbone_0.per_dout_val_1_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11492_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_2_ ),
    .Q(mem_backbone_0.per_dout_val_2_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11493_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_3_ ),
    .Q(mem_backbone_0.per_dout_val_3_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11494_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_4_ ),
    .Q(mem_backbone_0.per_dout_val_4_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11495_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_5_ ),
    .Q(mem_backbone_0.per_dout_val_5_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11496_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_6_ ),
    .Q(mem_backbone_0.per_dout_val_6_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11497_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_7_ ),
    .Q(mem_backbone_0.per_dout_val_7_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11498_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_8_ ),
    .Q(mem_backbone_0.per_dout_val_8_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11499_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_9_ ),
    .Q(mem_backbone_0.per_dout_val_9_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11500_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_10_ ),
    .Q(mem_backbone_0.per_dout_val_10_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11501_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_11_ ),
    .Q(mem_backbone_0.per_dout_val_11_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11502_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_12_ ),
    .Q(mem_backbone_0.per_dout_val_12_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11503_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_13_ ),
    .Q(mem_backbone_0.per_dout_val_13_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11504_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_14_ ),
    .Q(mem_backbone_0.per_dout_val_14_ ),
    .R(_04191_),
    .S(1'h1)
  );
  DFFSR _11505_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_15_ ),
    .Q(mem_backbone_0.per_dout_val_15_ ),
    .R(_04191_),
    .S(1'h1)
  );
  INVX1 _11506_ (
    .A(_00097_),
    .Y(_05103_)
  );
  INVX1 _11507_ (
    .A(_00104_),
    .Y(_05104_)
  );
  INVX1 _11508_ (
    .A(_00106_),
    .Y(_05105_)
  );
  INVX1 _11509_ (
    .A(_00107_),
    .Y(_05106_)
  );
  INVX1 _11510_ (
    .A(_00100_),
    .Y(_05107_)
  );
  INVX1 _11511_ (
    .A(multiplier_0.op2_0_ ),
    .Y(_05108_)
  );
  INVX1 _11512_ (
    .A(_00110_),
    .Y(_05109_)
  );
  INVX1 _11513_ (
    .A(multiplier_0.op2_1_ ),
    .Y(_05110_)
  );
  INVX1 _11514_ (
    .A(_00117_),
    .Y(_05111_)
  );
  INVX1 _11515_ (
    .A(multiplier_0.op2_2_ ),
    .Y(_05112_)
  );
  INVX1 _11516_ (
    .A(_00118_),
    .Y(_05113_)
  );
  INVX1 _11517_ (
    .A(multiplier_0.op2_3_ ),
    .Y(_05114_)
  );
  INVX1 _11518_ (
    .A(_00119_),
    .Y(_05115_)
  );
  INVX1 _11519_ (
    .A(multiplier_0.op2_4_ ),
    .Y(_05116_)
  );
  INVX1 _11520_ (
    .A(_00120_),
    .Y(_05117_)
  );
  INVX1 _11521_ (
    .A(multiplier_0.op2_5_ ),
    .Y(_05118_)
  );
  INVX1 _11522_ (
    .A(_00121_),
    .Y(_05119_)
  );
  INVX1 _11523_ (
    .A(multiplier_0.op2_6_ ),
    .Y(_05120_)
  );
  INVX1 _11524_ (
    .A(_00122_),
    .Y(_05121_)
  );
  INVX1 _11525_ (
    .A(multiplier_0.op2_7_ ),
    .Y(_05122_)
  );
  INVX1 _11526_ (
    .A(_00123_),
    .Y(_05123_)
  );
  INVX1 _11527_ (
    .A(multiplier_0.op1_0_ ),
    .Y(_05124_)
  );
  INVX1 _11528_ (
    .A(multiplier_0.op1_1_ ),
    .Y(_05125_)
  );
  INVX1 _11529_ (
    .A(multiplier_0.op1_2_ ),
    .Y(_05126_)
  );
  INVX1 _11530_ (
    .A(multiplier_0.op1_3_ ),
    .Y(_05127_)
  );
  INVX1 _11531_ (
    .A(multiplier_0.op1_4_ ),
    .Y(_05128_)
  );
  INVX1 _11532_ (
    .A(multiplier_0.op1_5_ ),
    .Y(_05129_)
  );
  INVX1 _11533_ (
    .A(multiplier_0.op1_6_ ),
    .Y(_05130_)
  );
  INVX1 _11534_ (
    .A(multiplier_0.op1_7_ ),
    .Y(_05131_)
  );
  INVX1 _11535_ (
    .A(multiplier_0.op1_8_ ),
    .Y(_05132_)
  );
  INVX1 _11536_ (
    .A(multiplier_0.op1_14_ ),
    .Y(_05133_)
  );
  INVX1 _11537_ (
    .A(multiplier_0.reslo_0_ ),
    .Y(_05134_)
  );
  INVX1 _11538_ (
    .A(multiplier_0.cycle_0_ ),
    .Y(_05135_)
  );
  INVX1 _11539_ (
    .A(multiplier_0.cycle_1_ ),
    .Y(_05136_)
  );
  INVX1 _11540_ (
    .A(multiplier_0.sign_sel ),
    .Y(_05137_)
  );
  INVX1 _11541_ (
    .A(multiplier_0.reslo_13_ ),
    .Y(_05138_)
  );
  INVX1 _11542_ (
    .A(multiplier_0.reslo_15_ ),
    .Y(_05139_)
  );
  INVX1 _11543_ (
    .A(multiplier_0.reshi_1_ ),
    .Y(_05140_)
  );
  INVX1 _11544_ (
    .A(multiplier_0.reshi_3_ ),
    .Y(_05141_)
  );
  INVX1 _11545_ (
    .A(multiplier_0.reshi_5_ ),
    .Y(_05142_)
  );
  INVX1 _11546_ (
    .A(multiplier_0.reshi_7_ ),
    .Y(_05143_)
  );
  INVX1 _11547_ (
    .A(multiplier_0.reshi_9_ ),
    .Y(_05144_)
  );
  INVX1 _11548_ (
    .A(multiplier_0.reshi_11_ ),
    .Y(_05145_)
  );
  INVX1 _11549_ (
    .A(multiplier_0.reshi_13_ ),
    .Y(_05146_)
  );
  INVX1 _11550_ (
    .A(_00162_),
    .Y(_04466_)
  );
  OR2X1 _11551_ (
    .A(_00099_),
    .B(1'h0),
    .Y(_05147_)
  );
  NAND2X1 _11552_ (
    .A(_05107_),
    .B(_00126_),
    .Y(_05148_)
  );
  NOR2X1 _11553_ (
    .A(_05147_),
    .B(_05148_),
    .Y(_05149_)
  );
  NOR2X1 _11554_ (
    .A(_00108_),
    .B(_05106_),
    .Y(_05150_)
  );
  NOR2X1 _11555_ (
    .A(_00098_),
    .B(_00109_),
    .Y(_05151_)
  );
  NAND2X1 _11556_ (
    .A(_05150_),
    .B(_05151_),
    .Y(_05152_)
  );
  NOR2X1 _11557_ (
    .A(_00106_),
    .B(_00105_),
    .Y(_05153_)
  );
  NAND3X1 _11558_ (
    .A(_00104_),
    .B(_00103_),
    .C(_05153_),
    .Y(_05154_)
  );
  NOR2X1 _11559_ (
    .A(_05152_),
    .B(_05154_),
    .Y(_05155_)
  );
  AND2X1 _11560_ (
    .A(_05149_),
    .B(_05155_),
    .Y(_05156_)
  );
  NOR2X1 _11561_ (
    .A(_00127_),
    .B(_00128_),
    .Y(_05157_)
  );
  OAI21X1 _11562_ (
    .A(_00127_),
    .B(_00128_),
    .C(_05156_),
    .Y(_05158_)
  );
  NAND2X1 _11563_ (
    .A(_05103_),
    .B(_00102_),
    .Y(_05159_)
  );
  OR2X1 _11564_ (
    .A(_00101_),
    .B(_05159_),
    .Y(_05160_)
  );
  OR2X1 _11565_ (
    .A(_05158_),
    .B(_05160_),
    .Y(_05161_)
  );
  INVX1 _11566_ (
    .A(_05161_),
    .Y(multiplier_0.op2_wr )
  );
  NOR2X1 _11567_ (
    .A(_05106_),
    .B(_00109_),
    .Y(_05162_)
  );
  NAND3X1 _11568_ (
    .A(_00103_),
    .B(_05105_),
    .C(_05162_),
    .Y(_05163_)
  );
  NOR2X1 _11569_ (
    .A(_00108_),
    .B(_00098_),
    .Y(_05164_)
  );
  NOR2X1 _11570_ (
    .A(_05104_),
    .B(_00105_),
    .Y(_05165_)
  );
  NAND3X1 _11571_ (
    .A(_05149_),
    .B(_05164_),
    .C(_05165_),
    .Y(_05166_)
  );
  NOR2X1 _11572_ (
    .A(_05163_),
    .B(_05166_),
    .Y(_05167_)
  );
  OAI21X1 _11573_ (
    .A(_00127_),
    .B(_00128_),
    .C(_05167_),
    .Y(_05168_)
  );
  OR2X1 _11574_ (
    .A(_05160_),
    .B(_05168_),
    .Y(_05169_)
  );
  MUX2X1 _11575_ (
    .A(multiplier_0.op2_0_ ),
    .B(_00110_),
    .S(_05169_),
    .Y(_05170_)
  );
  INVX1 _11576_ (
    .A(_05170_),
    .Y(_04415_)
  );
  MUX2X1 _11577_ (
    .A(multiplier_0.op2_1_ ),
    .B(_00117_),
    .S(_05169_),
    .Y(_05171_)
  );
  INVX1 _11578_ (
    .A(_05171_),
    .Y(_04422_)
  );
  MUX2X1 _11579_ (
    .A(multiplier_0.op2_2_ ),
    .B(_00118_),
    .S(_05169_),
    .Y(_05172_)
  );
  INVX1 _11580_ (
    .A(_05172_),
    .Y(_04423_)
  );
  MUX2X1 _11581_ (
    .A(multiplier_0.op2_3_ ),
    .B(_00119_),
    .S(_05169_),
    .Y(_05173_)
  );
  INVX1 _11582_ (
    .A(_05173_),
    .Y(_04424_)
  );
  MUX2X1 _11583_ (
    .A(multiplier_0.op2_4_ ),
    .B(_00120_),
    .S(_05169_),
    .Y(_05174_)
  );
  INVX1 _11584_ (
    .A(_05174_),
    .Y(_04425_)
  );
  MUX2X1 _11585_ (
    .A(multiplier_0.op2_5_ ),
    .B(_00121_),
    .S(_05169_),
    .Y(_05175_)
  );
  INVX1 _11586_ (
    .A(_05175_),
    .Y(_04426_)
  );
  MUX2X1 _11587_ (
    .A(multiplier_0.op2_6_ ),
    .B(_00122_),
    .S(_05169_),
    .Y(_05176_)
  );
  INVX1 _11588_ (
    .A(_05176_),
    .Y(_04427_)
  );
  MUX2X1 _11589_ (
    .A(multiplier_0.op2_7_ ),
    .B(_00123_),
    .S(_05169_),
    .Y(_05177_)
  );
  INVX1 _11590_ (
    .A(_05177_),
    .Y(_04428_)
  );
  OAI21X1 _11591_ (
    .A(_05158_),
    .B(_05160_),
    .C(multiplier_0.op2_8_ ),
    .Y(_05178_)
  );
  NAND2X1 _11592_ (
    .A(_00128_),
    .B(_00124_),
    .Y(_05179_)
  );
  OAI21X1 _11593_ (
    .A(_05169_),
    .B(_05179_),
    .C(_05178_),
    .Y(_04429_)
  );
  OAI21X1 _11594_ (
    .A(_05158_),
    .B(_05160_),
    .C(multiplier_0.op2_9_ ),
    .Y(_05180_)
  );
  NAND2X1 _11595_ (
    .A(_00128_),
    .B(_00125_),
    .Y(_05181_)
  );
  OAI21X1 _11596_ (
    .A(_05169_),
    .B(_05181_),
    .C(_05180_),
    .Y(_04430_)
  );
  OAI21X1 _11597_ (
    .A(_05158_),
    .B(_05160_),
    .C(multiplier_0.op2_10_ ),
    .Y(_05182_)
  );
  NAND2X1 _11598_ (
    .A(_00128_),
    .B(_00111_),
    .Y(_05183_)
  );
  OAI21X1 _11599_ (
    .A(_05169_),
    .B(_05183_),
    .C(_05182_),
    .Y(_04416_)
  );
  OAI21X1 _11600_ (
    .A(_05158_),
    .B(_05160_),
    .C(multiplier_0.op2_11_ ),
    .Y(_05184_)
  );
  NAND2X1 _11601_ (
    .A(_00128_),
    .B(_00112_),
    .Y(_05185_)
  );
  OAI21X1 _11602_ (
    .A(_05169_),
    .B(_05185_),
    .C(_05184_),
    .Y(_04417_)
  );
  OAI21X1 _11603_ (
    .A(_05158_),
    .B(_05160_),
    .C(multiplier_0.op2_12_ ),
    .Y(_05186_)
  );
  NAND2X1 _11604_ (
    .A(_00128_),
    .B(_00113_),
    .Y(_05187_)
  );
  OAI21X1 _11605_ (
    .A(_05169_),
    .B(_05187_),
    .C(_05186_),
    .Y(_04418_)
  );
  OAI21X1 _11606_ (
    .A(_05158_),
    .B(_05160_),
    .C(multiplier_0.op2_13_ ),
    .Y(_05188_)
  );
  NAND2X1 _11607_ (
    .A(_00128_),
    .B(_00114_),
    .Y(_05189_)
  );
  OAI21X1 _11608_ (
    .A(_05169_),
    .B(_05189_),
    .C(_05188_),
    .Y(_04419_)
  );
  OAI21X1 _11609_ (
    .A(_05158_),
    .B(_05160_),
    .C(multiplier_0.op2_14_ ),
    .Y(_05190_)
  );
  NAND2X1 _11610_ (
    .A(_00128_),
    .B(_00115_),
    .Y(_05191_)
  );
  OAI21X1 _11611_ (
    .A(_05169_),
    .B(_05191_),
    .C(_05190_),
    .Y(_04420_)
  );
  OAI21X1 _11612_ (
    .A(_05158_),
    .B(_05160_),
    .C(multiplier_0.op2_15_ ),
    .Y(_05192_)
  );
  NAND2X1 _11613_ (
    .A(_00128_),
    .B(_00116_),
    .Y(_05193_)
  );
  OAI21X1 _11614_ (
    .A(_05169_),
    .B(_05193_),
    .C(_05192_),
    .Y(_04421_)
  );
  OR2X1 _11615_ (
    .A(_00102_),
    .B(_05168_),
    .Y(_05194_)
  );
  MUX2X1 _11616_ (
    .A(multiplier_0.op1_0_ ),
    .B(_00110_),
    .S(_05194_),
    .Y(_05195_)
  );
  INVX1 _11617_ (
    .A(_05195_),
    .Y(_04399_)
  );
  MUX2X1 _11618_ (
    .A(multiplier_0.op1_1_ ),
    .B(_00117_),
    .S(_05194_),
    .Y(_05196_)
  );
  INVX1 _11619_ (
    .A(_05196_),
    .Y(_04406_)
  );
  MUX2X1 _11620_ (
    .A(multiplier_0.op1_2_ ),
    .B(_00118_),
    .S(_05194_),
    .Y(_05197_)
  );
  INVX1 _11621_ (
    .A(_05197_),
    .Y(_04407_)
  );
  MUX2X1 _11622_ (
    .A(multiplier_0.op1_3_ ),
    .B(_00119_),
    .S(_05194_),
    .Y(_05198_)
  );
  INVX1 _11623_ (
    .A(_05198_),
    .Y(_04408_)
  );
  MUX2X1 _11624_ (
    .A(multiplier_0.op1_4_ ),
    .B(_00120_),
    .S(_05194_),
    .Y(_05199_)
  );
  INVX1 _11625_ (
    .A(_05199_),
    .Y(_04409_)
  );
  MUX2X1 _11626_ (
    .A(multiplier_0.op1_5_ ),
    .B(_00121_),
    .S(_05194_),
    .Y(_05200_)
  );
  INVX1 _11627_ (
    .A(_05200_),
    .Y(_04410_)
  );
  MUX2X1 _11628_ (
    .A(multiplier_0.op1_6_ ),
    .B(_00122_),
    .S(_05194_),
    .Y(_05201_)
  );
  INVX1 _11629_ (
    .A(_05201_),
    .Y(_04411_)
  );
  MUX2X1 _11630_ (
    .A(multiplier_0.op1_7_ ),
    .B(_00123_),
    .S(_05194_),
    .Y(_05202_)
  );
  INVX1 _11631_ (
    .A(_05202_),
    .Y(_04412_)
  );
  OAI21X1 _11632_ (
    .A(_00102_),
    .B(_05158_),
    .C(multiplier_0.op1_8_ ),
    .Y(_05203_)
  );
  OAI21X1 _11633_ (
    .A(_05179_),
    .B(_05194_),
    .C(_05203_),
    .Y(_04413_)
  );
  OAI21X1 _11634_ (
    .A(_00102_),
    .B(_05158_),
    .C(multiplier_0.op1_9_ ),
    .Y(_05204_)
  );
  OAI21X1 _11635_ (
    .A(_05181_),
    .B(_05194_),
    .C(_05204_),
    .Y(_04414_)
  );
  OAI21X1 _11636_ (
    .A(_00102_),
    .B(_05158_),
    .C(multiplier_0.op1_10_ ),
    .Y(_05205_)
  );
  OAI21X1 _11637_ (
    .A(_05183_),
    .B(_05194_),
    .C(_05205_),
    .Y(_04400_)
  );
  OAI21X1 _11638_ (
    .A(_00102_),
    .B(_05158_),
    .C(multiplier_0.op1_11_ ),
    .Y(_05206_)
  );
  OAI21X1 _11639_ (
    .A(_05185_),
    .B(_05194_),
    .C(_05206_),
    .Y(_04401_)
  );
  OAI21X1 _11640_ (
    .A(_00102_),
    .B(_05158_),
    .C(multiplier_0.op1_12_ ),
    .Y(_05207_)
  );
  OAI21X1 _11641_ (
    .A(_05187_),
    .B(_05194_),
    .C(_05207_),
    .Y(_04402_)
  );
  OAI21X1 _11642_ (
    .A(_00102_),
    .B(_05158_),
    .C(multiplier_0.op1_13_ ),
    .Y(_05208_)
  );
  OAI21X1 _11643_ (
    .A(_05189_),
    .B(_05194_),
    .C(_05208_),
    .Y(_04403_)
  );
  OAI21X1 _11644_ (
    .A(_00102_),
    .B(_05158_),
    .C(multiplier_0.op1_14_ ),
    .Y(_05209_)
  );
  OAI21X1 _11645_ (
    .A(_05191_),
    .B(_05194_),
    .C(_05209_),
    .Y(_04404_)
  );
  OAI21X1 _11646_ (
    .A(_00102_),
    .B(_05158_),
    .C(multiplier_0.op1_15_ ),
    .Y(_05210_)
  );
  OAI21X1 _11647_ (
    .A(_05193_),
    .B(_05194_),
    .C(_05210_),
    .Y(_04405_)
  );
  NAND2X1 _11648_ (
    .A(multiplier_0.op2_8_ ),
    .B(multiplier_0.cycle_0_ ),
    .Y(_05211_)
  );
  OAI21X1 _11649_ (
    .A(_05108_),
    .B(multiplier_0.cycle_0_ ),
    .C(_05211_),
    .Y(_05212_)
  );
  MUX2X1 _11650_ (
    .A(multiplier_0.op2_8_ ),
    .B(multiplier_0.op2_0_ ),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05213_)
  );
  NAND3X1 _11651_ (
    .A(multiplier_0.op2_0_ ),
    .B(multiplier_0.op1_0_ ),
    .C(_05135_),
    .Y(_05214_)
  );
  NOR2X1 _11652_ (
    .A(_05136_),
    .B(_05214_),
    .Y(_05215_)
  );
  XNOR2X1 _11653_ (
    .A(_05134_),
    .B(_05215_),
    .Y(_05216_)
  );
  NAND2X1 _11654_ (
    .A(_00097_),
    .B(_00102_),
    .Y(_05217_)
  );
  OR2X1 _11655_ (
    .A(_00101_),
    .B(_05217_),
    .Y(_05218_)
  );
  OR2X1 _11656_ (
    .A(_05158_),
    .B(_05218_),
    .Y(_05219_)
  );
  INVX1 _11657_ (
    .A(_05219_),
    .Y(_05220_)
  );
  OAI21X1 _11658_ (
    .A(multiplier_0.acc_sel ),
    .B(_05161_),
    .C(_05219_),
    .Y(_05221_)
  );
  INVX1 _11659_ (
    .A(_05221_),
    .Y(_05222_)
  );
  NAND2X1 _11660_ (
    .A(_05216_),
    .B(_05222_),
    .Y(_05223_)
  );
  OAI21X1 _11661_ (
    .A(_05109_),
    .B(_05219_),
    .C(_05223_),
    .Y(_04447_)
  );
  NOR2X1 _11662_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.cycle_1_ ),
    .Y(_05224_)
  );
  NAND2X1 _11663_ (
    .A(_05135_),
    .B(_05136_),
    .Y(_05225_)
  );
  NOR2X1 _11664_ (
    .A(_05134_),
    .B(_05214_),
    .Y(_05226_)
  );
  INVX1 _11665_ (
    .A(_05226_),
    .Y(_05227_)
  );
  NAND2X1 _11666_ (
    .A(multiplier_0.op2_9_ ),
    .B(multiplier_0.cycle_0_ ),
    .Y(_05228_)
  );
  MUX2X1 _11667_ (
    .A(multiplier_0.op2_9_ ),
    .B(multiplier_0.op2_1_ ),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05229_)
  );
  OAI21X1 _11668_ (
    .A(_05110_),
    .B(multiplier_0.cycle_0_ ),
    .C(_05228_),
    .Y(_05230_)
  );
  OAI22X1 _11669_ (
    .A(_05125_),
    .B(_05213_),
    .C(_05229_),
    .D(_05124_),
    .Y(_05231_)
  );
  NOR2X1 _11670_ (
    .A(_05125_),
    .B(_05229_),
    .Y(_05232_)
  );
  NAND3X1 _11671_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05212_),
    .C(_05232_),
    .Y(_05233_)
  );
  NAND2X1 _11672_ (
    .A(_05231_),
    .B(_05233_),
    .Y(_05234_)
  );
  NOR2X1 _11673_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05234_),
    .Y(_05235_)
  );
  NAND2X1 _11674_ (
    .A(multiplier_0.reslo_1_ ),
    .B(_05235_),
    .Y(_05236_)
  );
  XNOR2X1 _11675_ (
    .A(multiplier_0.reslo_1_ ),
    .B(_05235_),
    .Y(_05237_)
  );
  XNOR2X1 _11676_ (
    .A(_05227_),
    .B(_05237_),
    .Y(_05238_)
  );
  OAI21X1 _11677_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.cycle_1_ ),
    .C(_05238_),
    .Y(_05239_)
  );
  OAI21X1 _11678_ (
    .A(multiplier_0.reslo_1_ ),
    .B(_05225_),
    .C(_05239_),
    .Y(_05240_)
  );
  NAND2X1 _11679_ (
    .A(_00117_),
    .B(_05220_),
    .Y(_05241_)
  );
  OAI21X1 _11680_ (
    .A(_05221_),
    .B(_05240_),
    .C(_05241_),
    .Y(_04454_)
  );
  OAI21X1 _11681_ (
    .A(_05227_),
    .B(_05237_),
    .C(_05236_),
    .Y(_05242_)
  );
  NAND2X1 _11682_ (
    .A(multiplier_0.op1_2_ ),
    .B(_05212_),
    .Y(_05243_)
  );
  NAND2X1 _11683_ (
    .A(multiplier_0.op2_10_ ),
    .B(multiplier_0.cycle_0_ ),
    .Y(_05244_)
  );
  MUX2X1 _11684_ (
    .A(multiplier_0.op2_10_ ),
    .B(multiplier_0.op2_2_ ),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05245_)
  );
  OAI21X1 _11685_ (
    .A(_05112_),
    .B(multiplier_0.cycle_0_ ),
    .C(_05244_),
    .Y(_05246_)
  );
  NOR2X1 _11686_ (
    .A(_05124_),
    .B(_05245_),
    .Y(_05247_)
  );
  NOR2X1 _11687_ (
    .A(_05125_),
    .B(_05245_),
    .Y(_05248_)
  );
  NAND2X1 _11688_ (
    .A(_05232_),
    .B(_05247_),
    .Y(_05249_)
  );
  XNOR2X1 _11689_ (
    .A(_05232_),
    .B(_05247_),
    .Y(_05250_)
  );
  XNOR2X1 _11690_ (
    .A(_05243_),
    .B(_05250_),
    .Y(_05251_)
  );
  NOR2X1 _11691_ (
    .A(_05233_),
    .B(_05251_),
    .Y(_05252_)
  );
  XNOR2X1 _11692_ (
    .A(_05233_),
    .B(_05251_),
    .Y(_05253_)
  );
  NOR2X1 _11693_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05253_),
    .Y(_05254_)
  );
  NAND2X1 _11694_ (
    .A(multiplier_0.reslo_2_ ),
    .B(_05254_),
    .Y(_05255_)
  );
  XOR2X1 _11695_ (
    .A(multiplier_0.reslo_2_ ),
    .B(_05254_),
    .Y(_05256_)
  );
  NAND2X1 _11696_ (
    .A(_05242_),
    .B(_05256_),
    .Y(_05257_)
  );
  XNOR2X1 _11697_ (
    .A(_05242_),
    .B(_05256_),
    .Y(_05258_)
  );
  OAI21X1 _11698_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.cycle_1_ ),
    .C(_05258_),
    .Y(_05259_)
  );
  OAI21X1 _11699_ (
    .A(multiplier_0.reslo_2_ ),
    .B(_05225_),
    .C(_05259_),
    .Y(_05260_)
  );
  NAND2X1 _11700_ (
    .A(_00118_),
    .B(_05220_),
    .Y(_05261_)
  );
  OAI21X1 _11701_ (
    .A(_05221_),
    .B(_05260_),
    .C(_05261_),
    .Y(_04455_)
  );
  NAND2X1 _11702_ (
    .A(_05255_),
    .B(_05257_),
    .Y(_05262_)
  );
  OAI21X1 _11703_ (
    .A(_05243_),
    .B(_05250_),
    .C(_05249_),
    .Y(_05263_)
  );
  INVX1 _11704_ (
    .A(_05263_),
    .Y(_05264_)
  );
  NAND2X1 _11705_ (
    .A(multiplier_0.op1_3_ ),
    .B(_05212_),
    .Y(_05265_)
  );
  NOR2X1 _11706_ (
    .A(_05126_),
    .B(_05229_),
    .Y(_05266_)
  );
  NOR2X1 _11707_ (
    .A(_05126_),
    .B(_05245_),
    .Y(_05267_)
  );
  NAND2X1 _11708_ (
    .A(_05232_),
    .B(_05267_),
    .Y(_05268_)
  );
  XNOR2X1 _11709_ (
    .A(_05248_),
    .B(_05266_),
    .Y(_05269_)
  );
  XNOR2X1 _11710_ (
    .A(_05265_),
    .B(_05269_),
    .Y(_05270_)
  );
  NOR2X1 _11711_ (
    .A(_05264_),
    .B(_05270_),
    .Y(_05271_)
  );
  INVX1 _11712_ (
    .A(_05271_),
    .Y(_05272_)
  );
  XOR2X1 _11713_ (
    .A(_05263_),
    .B(_05270_),
    .Y(_05273_)
  );
  NAND2X1 _11714_ (
    .A(multiplier_0.op2_11_ ),
    .B(multiplier_0.cycle_0_ ),
    .Y(_05274_)
  );
  MUX2X1 _11715_ (
    .A(multiplier_0.op2_11_ ),
    .B(multiplier_0.op2_3_ ),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05275_)
  );
  OAI21X1 _11716_ (
    .A(_05114_),
    .B(multiplier_0.cycle_0_ ),
    .C(_05274_),
    .Y(_05276_)
  );
  NAND2X1 _11717_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05276_),
    .Y(_05277_)
  );
  NOR2X1 _11718_ (
    .A(_05273_),
    .B(_05277_),
    .Y(_05278_)
  );
  XOR2X1 _11719_ (
    .A(_05273_),
    .B(_05277_),
    .Y(_05279_)
  );
  NAND2X1 _11720_ (
    .A(_05252_),
    .B(_05279_),
    .Y(_05280_)
  );
  XNOR2X1 _11721_ (
    .A(_05252_),
    .B(_05279_),
    .Y(_05281_)
  );
  NOR2X1 _11722_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05281_),
    .Y(_05282_)
  );
  AND2X1 _11723_ (
    .A(multiplier_0.reslo_3_ ),
    .B(_05282_),
    .Y(_05283_)
  );
  NOR2X1 _11724_ (
    .A(multiplier_0.reslo_3_ ),
    .B(_05282_),
    .Y(_05284_)
  );
  NOR2X1 _11725_ (
    .A(_05283_),
    .B(_05284_),
    .Y(_05285_)
  );
  XNOR2X1 _11726_ (
    .A(_05262_),
    .B(_05285_),
    .Y(_05286_)
  );
  OAI21X1 _11727_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.cycle_1_ ),
    .C(_05286_),
    .Y(_05287_)
  );
  OAI21X1 _11728_ (
    .A(multiplier_0.reslo_3_ ),
    .B(_05225_),
    .C(_05287_),
    .Y(_05288_)
  );
  NAND2X1 _11729_ (
    .A(_00119_),
    .B(_05220_),
    .Y(_05289_)
  );
  OAI21X1 _11730_ (
    .A(_05221_),
    .B(_05288_),
    .C(_05289_),
    .Y(_04456_)
  );
  AOI21X1 _11731_ (
    .A(_05262_),
    .B(_05285_),
    .C(_05283_),
    .Y(_05290_)
  );
  OAI21X1 _11732_ (
    .A(_05265_),
    .B(_05269_),
    .C(_05268_),
    .Y(_05291_)
  );
  NAND2X1 _11733_ (
    .A(multiplier_0.op1_4_ ),
    .B(_05212_),
    .Y(_05292_)
  );
  NOR2X1 _11734_ (
    .A(_05127_),
    .B(_05229_),
    .Y(_05293_)
  );
  NOR2X1 _11735_ (
    .A(_05127_),
    .B(_05245_),
    .Y(_05294_)
  );
  NAND2X1 _11736_ (
    .A(_05267_),
    .B(_05293_),
    .Y(_05295_)
  );
  XNOR2X1 _11737_ (
    .A(_05267_),
    .B(_05293_),
    .Y(_05296_)
  );
  XNOR2X1 _11738_ (
    .A(_05292_),
    .B(_05296_),
    .Y(_05297_)
  );
  INVX1 _11739_ (
    .A(_05297_),
    .Y(_05298_)
  );
  NAND2X1 _11740_ (
    .A(_05291_),
    .B(_05298_),
    .Y(_05299_)
  );
  XOR2X1 _11741_ (
    .A(_05291_),
    .B(_05297_),
    .Y(_05300_)
  );
  NAND2X1 _11742_ (
    .A(multiplier_0.op2_12_ ),
    .B(multiplier_0.cycle_0_ ),
    .Y(_05301_)
  );
  MUX2X1 _11743_ (
    .A(multiplier_0.op2_12_ ),
    .B(multiplier_0.op2_4_ ),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05302_)
  );
  OAI21X1 _11744_ (
    .A(_05116_),
    .B(multiplier_0.cycle_0_ ),
    .C(_05301_),
    .Y(_05303_)
  );
  NOR2X1 _11745_ (
    .A(_05125_),
    .B(_05302_),
    .Y(_05304_)
  );
  NAND3X1 _11746_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05276_),
    .C(_05304_),
    .Y(_05305_)
  );
  OAI22X1 _11747_ (
    .A(_05125_),
    .B(_05275_),
    .C(_05302_),
    .D(_05124_),
    .Y(_05306_)
  );
  NAND2X1 _11748_ (
    .A(_05305_),
    .B(_05306_),
    .Y(_05307_)
  );
  XOR2X1 _11749_ (
    .A(_05300_),
    .B(_05307_),
    .Y(_05308_)
  );
  NAND2X1 _11750_ (
    .A(_05278_),
    .B(_05308_),
    .Y(_05309_)
  );
  NOR2X1 _11751_ (
    .A(_05278_),
    .B(_05308_),
    .Y(_05310_)
  );
  XOR2X1 _11752_ (
    .A(_05278_),
    .B(_05308_),
    .Y(_05311_)
  );
  XNOR2X1 _11753_ (
    .A(_05271_),
    .B(_05311_),
    .Y(_05312_)
  );
  OR2X1 _11754_ (
    .A(_05280_),
    .B(_05312_),
    .Y(_05313_)
  );
  XOR2X1 _11755_ (
    .A(_05280_),
    .B(_05312_),
    .Y(_05314_)
  );
  NAND2X1 _11756_ (
    .A(_05135_),
    .B(_05314_),
    .Y(_05315_)
  );
  NAND3X1 _11757_ (
    .A(_05135_),
    .B(multiplier_0.reslo_4_ ),
    .C(_05314_),
    .Y(_05316_)
  );
  XOR2X1 _11758_ (
    .A(multiplier_0.reslo_4_ ),
    .B(_05315_),
    .Y(_05317_)
  );
  XNOR2X1 _11759_ (
    .A(_05290_),
    .B(_05317_),
    .Y(_05318_)
  );
  OAI21X1 _11760_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.cycle_1_ ),
    .C(_05318_),
    .Y(_05319_)
  );
  OAI21X1 _11761_ (
    .A(multiplier_0.reslo_4_ ),
    .B(_05225_),
    .C(_05319_),
    .Y(_05320_)
  );
  NAND2X1 _11762_ (
    .A(_00120_),
    .B(_05220_),
    .Y(_05321_)
  );
  OAI21X1 _11763_ (
    .A(_05221_),
    .B(_05320_),
    .C(_05321_),
    .Y(_04457_)
  );
  OAI21X1 _11764_ (
    .A(_05290_),
    .B(_05317_),
    .C(_05316_),
    .Y(_05322_)
  );
  OAI21X1 _11765_ (
    .A(_05272_),
    .B(_05310_),
    .C(_05309_),
    .Y(_05323_)
  );
  OAI21X1 _11766_ (
    .A(_05292_),
    .B(_05296_),
    .C(_05295_),
    .Y(_05324_)
  );
  NAND2X1 _11767_ (
    .A(multiplier_0.op1_5_ ),
    .B(_05212_),
    .Y(_05325_)
  );
  OR2X1 _11768_ (
    .A(_05128_),
    .B(_05229_),
    .Y(_05326_)
  );
  NAND3X1 _11769_ (
    .A(multiplier_0.op1_4_ ),
    .B(_05230_),
    .C(_05294_),
    .Y(_05327_)
  );
  XOR2X1 _11770_ (
    .A(_05294_),
    .B(_05326_),
    .Y(_05328_)
  );
  OR2X1 _11771_ (
    .A(_05325_),
    .B(_05328_),
    .Y(_05329_)
  );
  XNOR2X1 _11772_ (
    .A(_05325_),
    .B(_05328_),
    .Y(_05330_)
  );
  NOR2X1 _11773_ (
    .A(_05305_),
    .B(_05330_),
    .Y(_05331_)
  );
  XOR2X1 _11774_ (
    .A(_05305_),
    .B(_05330_),
    .Y(_05332_)
  );
  XNOR2X1 _11775_ (
    .A(_05324_),
    .B(_05332_),
    .Y(_05333_)
  );
  NAND2X1 _11776_ (
    .A(multiplier_0.op1_2_ ),
    .B(_05276_),
    .Y(_05334_)
  );
  NAND2X1 _11777_ (
    .A(multiplier_0.op2_13_ ),
    .B(multiplier_0.cycle_0_ ),
    .Y(_05335_)
  );
  MUX2X1 _11778_ (
    .A(multiplier_0.op2_13_ ),
    .B(multiplier_0.op2_5_ ),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05336_)
  );
  OAI21X1 _11779_ (
    .A(_05118_),
    .B(multiplier_0.cycle_0_ ),
    .C(_05335_),
    .Y(_05337_)
  );
  NOR2X1 _11780_ (
    .A(_05125_),
    .B(_05336_),
    .Y(_05338_)
  );
  NAND3X1 _11781_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05304_),
    .C(_05337_),
    .Y(_05339_)
  );
  AOI21X1 _11782_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05337_),
    .C(_05304_),
    .Y(_05340_)
  );
  OAI22X1 _11783_ (
    .A(_05125_),
    .B(_05302_),
    .C(_05336_),
    .D(_05124_),
    .Y(_05341_)
  );
  NAND2X1 _11784_ (
    .A(_05339_),
    .B(_05341_),
    .Y(_05342_)
  );
  XNOR2X1 _11785_ (
    .A(_05334_),
    .B(_05342_),
    .Y(_05343_)
  );
  NOR2X1 _11786_ (
    .A(_05333_),
    .B(_05343_),
    .Y(_05344_)
  );
  XOR2X1 _11787_ (
    .A(_05333_),
    .B(_05343_),
    .Y(_05345_)
  );
  OAI21X1 _11788_ (
    .A(_05300_),
    .B(_05307_),
    .C(_05299_),
    .Y(_05346_)
  );
  NAND2X1 _11789_ (
    .A(_05345_),
    .B(_05346_),
    .Y(_05347_)
  );
  XOR2X1 _11790_ (
    .A(_05345_),
    .B(_05346_),
    .Y(_05348_)
  );
  NAND2X1 _11791_ (
    .A(_05323_),
    .B(_05348_),
    .Y(_05349_)
  );
  INVX1 _11792_ (
    .A(_05349_),
    .Y(_05350_)
  );
  XNOR2X1 _11793_ (
    .A(_05323_),
    .B(_05348_),
    .Y(_05351_)
  );
  NOR2X1 _11794_ (
    .A(_05313_),
    .B(_05351_),
    .Y(_05352_)
  );
  XNOR2X1 _11795_ (
    .A(_05313_),
    .B(_05351_),
    .Y(_05353_)
  );
  NOR2X1 _11796_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05353_),
    .Y(_05354_)
  );
  AND2X1 _11797_ (
    .A(multiplier_0.reslo_5_ ),
    .B(_05354_),
    .Y(_05355_)
  );
  XOR2X1 _11798_ (
    .A(multiplier_0.reslo_5_ ),
    .B(_05354_),
    .Y(_05356_)
  );
  XNOR2X1 _11799_ (
    .A(_05322_),
    .B(_05356_),
    .Y(_05357_)
  );
  OAI21X1 _11800_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.cycle_1_ ),
    .C(_05357_),
    .Y(_05358_)
  );
  OAI21X1 _11801_ (
    .A(multiplier_0.reslo_5_ ),
    .B(_05225_),
    .C(_05358_),
    .Y(_05359_)
  );
  NAND2X1 _11802_ (
    .A(_00121_),
    .B(_05220_),
    .Y(_05360_)
  );
  OAI21X1 _11803_ (
    .A(_05221_),
    .B(_05359_),
    .C(_05360_),
    .Y(_04458_)
  );
  AOI21X1 _11804_ (
    .A(_05322_),
    .B(_05356_),
    .C(_05355_),
    .Y(_05361_)
  );
  AOI21X1 _11805_ (
    .A(_05324_),
    .B(_05332_),
    .C(_05331_),
    .Y(_05362_)
  );
  OAI21X1 _11806_ (
    .A(_05325_),
    .B(_05328_),
    .C(_05327_),
    .Y(_05363_)
  );
  NAND2X1 _11807_ (
    .A(multiplier_0.op1_6_ ),
    .B(_05212_),
    .Y(_05364_)
  );
  NOR2X1 _11808_ (
    .A(_05129_),
    .B(_05245_),
    .Y(_05365_)
  );
  OR2X1 _11809_ (
    .A(_05129_),
    .B(_05245_),
    .Y(_05366_)
  );
  OAI22X1 _11810_ (
    .A(_05129_),
    .B(_05229_),
    .C(_05245_),
    .D(_05128_),
    .Y(_05367_)
  );
  OAI21X1 _11811_ (
    .A(_05326_),
    .B(_05366_),
    .C(_05367_),
    .Y(_05368_)
  );
  XNOR2X1 _11812_ (
    .A(_05364_),
    .B(_05368_),
    .Y(_05369_)
  );
  OAI21X1 _11813_ (
    .A(_05334_),
    .B(_05340_),
    .C(_05339_),
    .Y(_05370_)
  );
  INVX1 _11814_ (
    .A(_05370_),
    .Y(_05371_)
  );
  NOR2X1 _11815_ (
    .A(_05369_),
    .B(_05371_),
    .Y(_05372_)
  );
  XOR2X1 _11816_ (
    .A(_05369_),
    .B(_05370_),
    .Y(_05373_)
  );
  AOI21X1 _11817_ (
    .A(_05327_),
    .B(_05329_),
    .C(_05373_),
    .Y(_05374_)
  );
  XOR2X1 _11818_ (
    .A(_05363_),
    .B(_05373_),
    .Y(_05375_)
  );
  NAND2X1 _11819_ (
    .A(multiplier_0.op1_3_ ),
    .B(_05276_),
    .Y(_05376_)
  );
  NOR2X1 _11820_ (
    .A(_05126_),
    .B(_05302_),
    .Y(_05377_)
  );
  NOR2X1 _11821_ (
    .A(_05126_),
    .B(_05336_),
    .Y(_05378_)
  );
  NAND2X1 _11822_ (
    .A(_05304_),
    .B(_05378_),
    .Y(_05379_)
  );
  XNOR2X1 _11823_ (
    .A(_05338_),
    .B(_05377_),
    .Y(_05380_)
  );
  XNOR2X1 _11824_ (
    .A(_05376_),
    .B(_05380_),
    .Y(_05381_)
  );
  NAND2X1 _11825_ (
    .A(multiplier_0.op2_14_ ),
    .B(multiplier_0.cycle_0_ ),
    .Y(_05382_)
  );
  MUX2X1 _11826_ (
    .A(multiplier_0.op2_14_ ),
    .B(multiplier_0.op2_6_ ),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05383_)
  );
  OAI21X1 _11827_ (
    .A(_05120_),
    .B(multiplier_0.cycle_0_ ),
    .C(_05382_),
    .Y(_05384_)
  );
  NAND2X1 _11828_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05384_),
    .Y(_05385_)
  );
  NOR2X1 _11829_ (
    .A(_05381_),
    .B(_05385_),
    .Y(_05386_)
  );
  XNOR2X1 _11830_ (
    .A(_05381_),
    .B(_05385_),
    .Y(_05387_)
  );
  NOR2X1 _11831_ (
    .A(_05375_),
    .B(_05387_),
    .Y(_05388_)
  );
  XOR2X1 _11832_ (
    .A(_05375_),
    .B(_05387_),
    .Y(_05389_)
  );
  NAND2X1 _11833_ (
    .A(_05344_),
    .B(_05389_),
    .Y(_05390_)
  );
  XNOR2X1 _11834_ (
    .A(_05344_),
    .B(_05389_),
    .Y(_05391_)
  );
  XOR2X1 _11835_ (
    .A(_05362_),
    .B(_05391_),
    .Y(_05392_)
  );
  NAND3X1 _11836_ (
    .A(_05345_),
    .B(_05346_),
    .C(_05392_),
    .Y(_05393_)
  );
  XNOR2X1 _11837_ (
    .A(_05347_),
    .B(_05392_),
    .Y(_05394_)
  );
  XNOR2X1 _11838_ (
    .A(_05352_),
    .B(_05394_),
    .Y(_05395_)
  );
  MUX2X1 _11839_ (
    .A(_05394_),
    .B(_05395_),
    .S(_05350_),
    .Y(_05396_)
  );
  NAND2X1 _11840_ (
    .A(_05135_),
    .B(_05396_),
    .Y(_05397_)
  );
  NAND3X1 _11841_ (
    .A(_05135_),
    .B(multiplier_0.reslo_6_ ),
    .C(_05396_),
    .Y(_05398_)
  );
  AOI21X1 _11842_ (
    .A(_05135_),
    .B(_05396_),
    .C(multiplier_0.reslo_6_ ),
    .Y(_05399_)
  );
  XNOR2X1 _11843_ (
    .A(multiplier_0.reslo_6_ ),
    .B(_05397_),
    .Y(_05400_)
  );
  XOR2X1 _11844_ (
    .A(_05361_),
    .B(_05400_),
    .Y(_05401_)
  );
  OAI21X1 _11845_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.cycle_1_ ),
    .C(_05401_),
    .Y(_05402_)
  );
  OAI21X1 _11846_ (
    .A(multiplier_0.reslo_6_ ),
    .B(_05225_),
    .C(_05402_),
    .Y(_05403_)
  );
  NAND2X1 _11847_ (
    .A(_00122_),
    .B(_05220_),
    .Y(_05404_)
  );
  OAI21X1 _11848_ (
    .A(_05221_),
    .B(_05403_),
    .C(_05404_),
    .Y(_04459_)
  );
  OAI21X1 _11849_ (
    .A(_05361_),
    .B(_05399_),
    .C(_05398_),
    .Y(_05405_)
  );
  OAI21X1 _11850_ (
    .A(_05350_),
    .B(_05352_),
    .C(_05394_),
    .Y(_05406_)
  );
  OAI21X1 _11851_ (
    .A(_05362_),
    .B(_05391_),
    .C(_05390_),
    .Y(_05407_)
  );
  NOR2X1 _11852_ (
    .A(_05372_),
    .B(_05374_),
    .Y(_05408_)
  );
  OAI22X1 _11853_ (
    .A(_05326_),
    .B(_05366_),
    .C(_05368_),
    .D(_05364_),
    .Y(_05409_)
  );
  NAND2X1 _11854_ (
    .A(multiplier_0.op1_7_ ),
    .B(_05212_),
    .Y(_05410_)
  );
  NOR2X1 _11855_ (
    .A(_05130_),
    .B(_05229_),
    .Y(_05411_)
  );
  NAND2X1 _11856_ (
    .A(_05365_),
    .B(_05411_),
    .Y(_05412_)
  );
  XNOR2X1 _11857_ (
    .A(_05365_),
    .B(_05411_),
    .Y(_05413_)
  );
  XNOR2X1 _11858_ (
    .A(_05410_),
    .B(_05413_),
    .Y(_05414_)
  );
  INVX1 _11859_ (
    .A(_05414_),
    .Y(_05415_)
  );
  OAI21X1 _11860_ (
    .A(_05376_),
    .B(_05380_),
    .C(_05379_),
    .Y(_05416_)
  );
  NAND2X1 _11861_ (
    .A(_05415_),
    .B(_05416_),
    .Y(_05417_)
  );
  XOR2X1 _11862_ (
    .A(_05414_),
    .B(_05416_),
    .Y(_05418_)
  );
  INVX1 _11863_ (
    .A(_05418_),
    .Y(_05419_)
  );
  NAND2X1 _11864_ (
    .A(_05409_),
    .B(_05419_),
    .Y(_05420_)
  );
  XOR2X1 _11865_ (
    .A(_05409_),
    .B(_05418_),
    .Y(_05421_)
  );
  NAND2X1 _11866_ (
    .A(multiplier_0.op1_4_ ),
    .B(_05276_),
    .Y(_05422_)
  );
  NOR2X1 _11867_ (
    .A(_05127_),
    .B(_05302_),
    .Y(_05423_)
  );
  NOR2X1 _11868_ (
    .A(_05127_),
    .B(_05336_),
    .Y(_05424_)
  );
  NAND2X1 _11869_ (
    .A(_05377_),
    .B(_05424_),
    .Y(_05425_)
  );
  XNOR2X1 _11870_ (
    .A(_05378_),
    .B(_05423_),
    .Y(_05426_)
  );
  XNOR2X1 _11871_ (
    .A(_05422_),
    .B(_05426_),
    .Y(_05427_)
  );
  NAND2X1 _11872_ (
    .A(multiplier_0.op2_15_ ),
    .B(multiplier_0.cycle_0_ ),
    .Y(_05428_)
  );
  MUX2X1 _11873_ (
    .A(multiplier_0.op2_15_ ),
    .B(multiplier_0.op2_7_ ),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05429_)
  );
  OAI21X1 _11874_ (
    .A(_05122_),
    .B(multiplier_0.cycle_0_ ),
    .C(_05428_),
    .Y(_05430_)
  );
  OAI22X1 _11875_ (
    .A(_05125_),
    .B(_05383_),
    .C(_05429_),
    .D(_05124_),
    .Y(_05431_)
  );
  NOR2X1 _11876_ (
    .A(_05125_),
    .B(_05429_),
    .Y(_05432_)
  );
  NAND3X1 _11877_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05384_),
    .C(_05432_),
    .Y(_05433_)
  );
  NAND2X1 _11878_ (
    .A(_05431_),
    .B(_05433_),
    .Y(_05434_)
  );
  NOR2X1 _11879_ (
    .A(_05427_),
    .B(_05434_),
    .Y(_05435_)
  );
  XOR2X1 _11880_ (
    .A(_05427_),
    .B(_05434_),
    .Y(_05436_)
  );
  NAND2X1 _11881_ (
    .A(_05386_),
    .B(_05436_),
    .Y(_05437_)
  );
  XNOR2X1 _11882_ (
    .A(_05386_),
    .B(_05436_),
    .Y(_05438_)
  );
  XOR2X1 _11883_ (
    .A(_05421_),
    .B(_05438_),
    .Y(_05439_)
  );
  NAND2X1 _11884_ (
    .A(_05388_),
    .B(_05439_),
    .Y(_05440_)
  );
  XNOR2X1 _11885_ (
    .A(_05388_),
    .B(_05439_),
    .Y(_05441_)
  );
  XOR2X1 _11886_ (
    .A(_05408_),
    .B(_05441_),
    .Y(_05442_)
  );
  NAND2X1 _11887_ (
    .A(_05407_),
    .B(_05442_),
    .Y(_05443_)
  );
  XNOR2X1 _11888_ (
    .A(_05407_),
    .B(_05442_),
    .Y(_05444_)
  );
  OR2X1 _11889_ (
    .A(_05393_),
    .B(_05444_),
    .Y(_05445_)
  );
  AND2X1 _11890_ (
    .A(_05393_),
    .B(_05444_),
    .Y(_05446_)
  );
  XNOR2X1 _11891_ (
    .A(_05393_),
    .B(_05444_),
    .Y(_05447_)
  );
  XNOR2X1 _11892_ (
    .A(_05406_),
    .B(_05447_),
    .Y(_05448_)
  );
  NOR2X1 _11893_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05448_),
    .Y(_05449_)
  );
  AND2X1 _11894_ (
    .A(multiplier_0.reslo_7_ ),
    .B(_05449_),
    .Y(_05450_)
  );
  XOR2X1 _11895_ (
    .A(multiplier_0.reslo_7_ ),
    .B(_05449_),
    .Y(_05451_)
  );
  XNOR2X1 _11896_ (
    .A(_05405_),
    .B(_05451_),
    .Y(_05452_)
  );
  OAI21X1 _11897_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.cycle_1_ ),
    .C(_05452_),
    .Y(_05453_)
  );
  OAI21X1 _11898_ (
    .A(multiplier_0.reslo_7_ ),
    .B(_05225_),
    .C(_05453_),
    .Y(_05454_)
  );
  NAND2X1 _11899_ (
    .A(_00123_),
    .B(_05220_),
    .Y(_05455_)
  );
  OAI21X1 _11900_ (
    .A(_05221_),
    .B(_05454_),
    .C(_05455_),
    .Y(_04460_)
  );
  AOI21X1 _11901_ (
    .A(_05405_),
    .B(_05451_),
    .C(_05450_),
    .Y(_05456_)
  );
  OR2X1 _11902_ (
    .A(_05124_),
    .B(_05211_),
    .Y(_05457_)
  );
  OAI21X1 _11903_ (
    .A(_05406_),
    .B(_05446_),
    .C(_05445_),
    .Y(_05458_)
  );
  NAND2X1 _11904_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05212_),
    .Y(_05459_)
  );
  OAI21X1 _11905_ (
    .A(_05408_),
    .B(_05441_),
    .C(_05440_),
    .Y(_05460_)
  );
  NAND2X1 _11906_ (
    .A(_05417_),
    .B(_05420_),
    .Y(_05461_)
  );
  OAI21X1 _11907_ (
    .A(_05421_),
    .B(_05438_),
    .C(_05437_),
    .Y(_05462_)
  );
  OAI21X1 _11908_ (
    .A(_05410_),
    .B(_05413_),
    .C(_05412_),
    .Y(_05463_)
  );
  INVX1 _11909_ (
    .A(_05463_),
    .Y(_05464_)
  );
  NAND2X1 _11910_ (
    .A(multiplier_0.op1_7_ ),
    .B(_05230_),
    .Y(_05465_)
  );
  OR2X1 _11911_ (
    .A(_05130_),
    .B(_05275_),
    .Y(_05466_)
  );
  OAI22X1 _11912_ (
    .A(_05130_),
    .B(_05245_),
    .C(_05275_),
    .D(_05129_),
    .Y(_05467_)
  );
  OAI21X1 _11913_ (
    .A(_05366_),
    .B(_05466_),
    .C(_05467_),
    .Y(_05468_)
  );
  XNOR2X1 _11914_ (
    .A(_05465_),
    .B(_05468_),
    .Y(_05469_)
  );
  INVX1 _11915_ (
    .A(_05469_),
    .Y(_05470_)
  );
  OAI21X1 _11916_ (
    .A(_05422_),
    .B(_05426_),
    .C(_05425_),
    .Y(_05471_)
  );
  NAND2X1 _11917_ (
    .A(_05470_),
    .B(_05471_),
    .Y(_05472_)
  );
  XOR2X1 _11918_ (
    .A(_05469_),
    .B(_05471_),
    .Y(_05473_)
  );
  XNOR2X1 _11919_ (
    .A(_05464_),
    .B(_05473_),
    .Y(_05474_)
  );
  NAND2X1 _11920_ (
    .A(multiplier_0.op1_4_ ),
    .B(_05303_),
    .Y(_05475_)
  );
  NOR2X1 _11921_ (
    .A(_05126_),
    .B(_05383_),
    .Y(_05476_)
  );
  NAND2X1 _11922_ (
    .A(multiplier_0.op1_3_ ),
    .B(_05384_),
    .Y(_05477_)
  );
  NAND2X1 _11923_ (
    .A(_05424_),
    .B(_05476_),
    .Y(_05478_)
  );
  XNOR2X1 _11924_ (
    .A(_05424_),
    .B(_05476_),
    .Y(_05479_)
  );
  XNOR2X1 _11925_ (
    .A(_05475_),
    .B(_05479_),
    .Y(_05480_)
  );
  NAND3X1 _11926_ (
    .A(multiplier_0.op2_15_ ),
    .B(multiplier_0.cycle_0_ ),
    .C(multiplier_0.sign_sel ),
    .Y(_05481_)
  );
  INVX1 _11927_ (
    .A(_05481_),
    .Y(_05482_)
  );
  NAND2X1 _11928_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05482_),
    .Y(_05483_)
  );
  OAI21X1 _11929_ (
    .A(_05124_),
    .B(_05383_),
    .C(_05432_),
    .Y(_05484_)
  );
  XNOR2X1 _11930_ (
    .A(_05483_),
    .B(_05484_),
    .Y(_05485_)
  );
  XOR2X1 _11931_ (
    .A(_05480_),
    .B(_05485_),
    .Y(_05486_)
  );
  NAND2X1 _11932_ (
    .A(_05435_),
    .B(_05486_),
    .Y(_05487_)
  );
  XNOR2X1 _11933_ (
    .A(_05435_),
    .B(_05486_),
    .Y(_05488_)
  );
  XOR2X1 _11934_ (
    .A(_05474_),
    .B(_05488_),
    .Y(_05489_)
  );
  AND2X1 _11935_ (
    .A(_05462_),
    .B(_05489_),
    .Y(_05490_)
  );
  XNOR2X1 _11936_ (
    .A(_05462_),
    .B(_05489_),
    .Y(_05491_)
  );
  AOI21X1 _11937_ (
    .A(_05417_),
    .B(_05420_),
    .C(_05491_),
    .Y(_05492_)
  );
  XOR2X1 _11938_ (
    .A(_05461_),
    .B(_05491_),
    .Y(_05493_)
  );
  INVX1 _11939_ (
    .A(_05493_),
    .Y(_05494_)
  );
  AND2X1 _11940_ (
    .A(_05460_),
    .B(_05494_),
    .Y(_05495_)
  );
  NAND2X1 _11941_ (
    .A(_05460_),
    .B(_05494_),
    .Y(_05496_)
  );
  XOR2X1 _11942_ (
    .A(_05460_),
    .B(_05493_),
    .Y(_05497_)
  );
  NOR2X1 _11943_ (
    .A(_05459_),
    .B(_05497_),
    .Y(_05498_)
  );
  OR2X1 _11944_ (
    .A(_05459_),
    .B(_05497_),
    .Y(_05499_)
  );
  XNOR2X1 _11945_ (
    .A(_05459_),
    .B(_05497_),
    .Y(_05500_)
  );
  NOR2X1 _11946_ (
    .A(_05443_),
    .B(_05500_),
    .Y(_05501_)
  );
  XOR2X1 _11947_ (
    .A(_05443_),
    .B(_05500_),
    .Y(_05502_)
  );
  XNOR2X1 _11948_ (
    .A(_05458_),
    .B(_05502_),
    .Y(_05503_)
  );
  OAI21X1 _11949_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05503_),
    .C(_05457_),
    .Y(_05504_)
  );
  NAND2X1 _11950_ (
    .A(multiplier_0.reslo_8_ ),
    .B(_05504_),
    .Y(_05505_)
  );
  XNOR2X1 _11951_ (
    .A(multiplier_0.reslo_8_ ),
    .B(_05504_),
    .Y(_05506_)
  );
  XOR2X1 _11952_ (
    .A(_05456_),
    .B(_05506_),
    .Y(_05507_)
  );
  NOR2X1 _11953_ (
    .A(_05224_),
    .B(_05507_),
    .Y(_05508_)
  );
  OAI21X1 _11954_ (
    .A(multiplier_0.reslo_8_ ),
    .B(_05225_),
    .C(_05222_),
    .Y(_05509_)
  );
  OAI22X1 _11955_ (
    .A(_05179_),
    .B(_05219_),
    .C(_05508_),
    .D(_05509_),
    .Y(_04461_)
  );
  OAI21X1 _11956_ (
    .A(_05456_),
    .B(_05506_),
    .C(_05505_),
    .Y(_05510_)
  );
  AOI21X1 _11957_ (
    .A(_05458_),
    .B(_05502_),
    .C(_05501_),
    .Y(_05511_)
  );
  OR2X1 _11958_ (
    .A(_05490_),
    .B(_05492_),
    .Y(_05512_)
  );
  OAI21X1 _11959_ (
    .A(_05464_),
    .B(_05473_),
    .C(_05472_),
    .Y(_05513_)
  );
  INVX1 _11960_ (
    .A(_05513_),
    .Y(_05514_)
  );
  OAI21X1 _11961_ (
    .A(_05474_),
    .B(_05488_),
    .C(_05487_),
    .Y(_05515_)
  );
  OAI22X1 _11962_ (
    .A(_05366_),
    .B(_05466_),
    .C(_05468_),
    .D(_05465_),
    .Y(_05516_)
  );
  NAND2X1 _11963_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05212_),
    .Y(_05517_)
  );
  OAI22X1 _11964_ (
    .A(_05132_),
    .B(_05229_),
    .C(_05245_),
    .D(_05131_),
    .Y(_05518_)
  );
  NAND2X1 _11965_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05246_),
    .Y(_05519_)
  );
  NOR2X1 _11966_ (
    .A(_05465_),
    .B(_05519_),
    .Y(_05520_)
  );
  OAI21X1 _11967_ (
    .A(_05465_),
    .B(_05519_),
    .C(_05518_),
    .Y(_05521_)
  );
  NOR2X1 _11968_ (
    .A(_05517_),
    .B(_05521_),
    .Y(_05522_)
  );
  XNOR2X1 _11969_ (
    .A(_05517_),
    .B(_05521_),
    .Y(_05523_)
  );
  INVX1 _11970_ (
    .A(_05523_),
    .Y(_05524_)
  );
  OAI21X1 _11971_ (
    .A(_05475_),
    .B(_05479_),
    .C(_05478_),
    .Y(_05525_)
  );
  NAND2X1 _11972_ (
    .A(_05524_),
    .B(_05525_),
    .Y(_05526_)
  );
  XOR2X1 _11973_ (
    .A(_05523_),
    .B(_05525_),
    .Y(_05527_)
  );
  INVX1 _11974_ (
    .A(_05527_),
    .Y(_05528_)
  );
  NAND2X1 _11975_ (
    .A(_05516_),
    .B(_05528_),
    .Y(_05529_)
  );
  XOR2X1 _11976_ (
    .A(_05516_),
    .B(_05527_),
    .Y(_05530_)
  );
  OAI22X1 _11977_ (
    .A(_05433_),
    .B(_05482_),
    .C(_05485_),
    .D(_05480_),
    .Y(_05531_)
  );
  NAND2X1 _11978_ (
    .A(multiplier_0.op1_5_ ),
    .B(_05337_),
    .Y(_05532_)
  );
  OAI22X1 _11979_ (
    .A(_05129_),
    .B(_05302_),
    .C(_05336_),
    .D(_05128_),
    .Y(_05533_)
  );
  OAI21X1 _11980_ (
    .A(_05475_),
    .B(_05532_),
    .C(_05533_),
    .Y(_05534_)
  );
  XNOR2X1 _11981_ (
    .A(_05466_),
    .B(_05534_),
    .Y(_05535_)
  );
  INVX1 _11982_ (
    .A(_05535_),
    .Y(_05536_)
  );
  OAI21X1 _11983_ (
    .A(_05124_),
    .B(_05432_),
    .C(_05482_),
    .Y(_05537_)
  );
  NOR2X1 _11984_ (
    .A(_05126_),
    .B(_05429_),
    .Y(_05538_)
  );
  NOR2X1 _11985_ (
    .A(multiplier_0.op1_1_ ),
    .B(_05481_),
    .Y(_05539_)
  );
  XNOR2X1 _11986_ (
    .A(_05538_),
    .B(_05539_),
    .Y(_05540_)
  );
  NOR2X1 _11987_ (
    .A(_05477_),
    .B(_05540_),
    .Y(_05541_)
  );
  XNOR2X1 _11988_ (
    .A(_05477_),
    .B(_05540_),
    .Y(_05542_)
  );
  XOR2X1 _11989_ (
    .A(_05537_),
    .B(_05542_),
    .Y(_05543_)
  );
  NAND2X1 _11990_ (
    .A(_05536_),
    .B(_05543_),
    .Y(_05544_)
  );
  XNOR2X1 _11991_ (
    .A(_05535_),
    .B(_05543_),
    .Y(_05545_)
  );
  NAND2X1 _11992_ (
    .A(_05531_),
    .B(_05545_),
    .Y(_05546_)
  );
  XNOR2X1 _11993_ (
    .A(_05531_),
    .B(_05545_),
    .Y(_05547_)
  );
  XOR2X1 _11994_ (
    .A(_05530_),
    .B(_05547_),
    .Y(_05548_)
  );
  NAND2X1 _11995_ (
    .A(_05515_),
    .B(_05548_),
    .Y(_05549_)
  );
  XNOR2X1 _11996_ (
    .A(_05515_),
    .B(_05548_),
    .Y(_05550_)
  );
  XNOR2X1 _11997_ (
    .A(_05514_),
    .B(_05550_),
    .Y(_05551_)
  );
  INVX1 _11998_ (
    .A(_05551_),
    .Y(_05552_)
  );
  OAI21X1 _11999_ (
    .A(_05490_),
    .B(_05492_),
    .C(_05552_),
    .Y(_05553_)
  );
  XNOR2X1 _12000_ (
    .A(_05512_),
    .B(_05551_),
    .Y(_05554_)
  );
  XOR2X1 _12001_ (
    .A(_05512_),
    .B(_05551_),
    .Y(_05555_)
  );
  OAI21X1 _12002_ (
    .A(_05495_),
    .B(_05498_),
    .C(_05554_),
    .Y(_05556_)
  );
  NAND3X1 _12003_ (
    .A(_05496_),
    .B(_05499_),
    .C(_05555_),
    .Y(_05557_)
  );
  INVX1 _12004_ (
    .A(_05557_),
    .Y(_05558_)
  );
  NAND2X1 _12005_ (
    .A(_05556_),
    .B(_05557_),
    .Y(_05559_)
  );
  XNOR2X1 _12006_ (
    .A(_05511_),
    .B(_05559_),
    .Y(_05560_)
  );
  MUX2X1 _12007_ (
    .A(_05234_),
    .B(_05560_),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05561_)
  );
  OR2X1 _12008_ (
    .A(multiplier_0.reslo_9_ ),
    .B(_05561_),
    .Y(_05562_)
  );
  AND2X1 _12009_ (
    .A(multiplier_0.reslo_9_ ),
    .B(_05561_),
    .Y(_05563_)
  );
  NAND2X1 _12010_ (
    .A(multiplier_0.reslo_9_ ),
    .B(_05561_),
    .Y(_05564_)
  );
  NAND2X1 _12011_ (
    .A(_05562_),
    .B(_05564_),
    .Y(_05565_)
  );
  XNOR2X1 _12012_ (
    .A(_05510_),
    .B(_05565_),
    .Y(_05566_)
  );
  NOR2X1 _12013_ (
    .A(_05224_),
    .B(_05566_),
    .Y(_05567_)
  );
  OAI21X1 _12014_ (
    .A(multiplier_0.reslo_9_ ),
    .B(_05225_),
    .C(_05222_),
    .Y(_05568_)
  );
  OAI22X1 _12015_ (
    .A(_05181_),
    .B(_05219_),
    .C(_05567_),
    .D(_05568_),
    .Y(_04462_)
  );
  AOI21X1 _12016_ (
    .A(_05510_),
    .B(_05562_),
    .C(_05563_),
    .Y(_05569_)
  );
  OAI21X1 _12017_ (
    .A(_05514_),
    .B(_05550_),
    .C(_05549_),
    .Y(_05570_)
  );
  NAND2X1 _12018_ (
    .A(_05526_),
    .B(_05529_),
    .Y(_05571_)
  );
  OAI21X1 _12019_ (
    .A(_05530_),
    .B(_05547_),
    .C(_05546_),
    .Y(_05572_)
  );
  INVX1 _12020_ (
    .A(_05572_),
    .Y(_05573_)
  );
  NOR2X1 _12021_ (
    .A(_05520_),
    .B(_05522_),
    .Y(_05574_)
  );
  NAND2X1 _12022_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05212_),
    .Y(_05575_)
  );
  NAND2X1 _12023_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05230_),
    .Y(_05576_)
  );
  AND2X1 _12024_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05246_),
    .Y(_05577_)
  );
  OR2X1 _12025_ (
    .A(_05519_),
    .B(_05576_),
    .Y(_05578_)
  );
  XNOR2X1 _12026_ (
    .A(_05519_),
    .B(_05576_),
    .Y(_05579_)
  );
  OR2X1 _12027_ (
    .A(_05575_),
    .B(_05579_),
    .Y(_05580_)
  );
  NAND2X1 _12028_ (
    .A(_05575_),
    .B(_05579_),
    .Y(_05581_)
  );
  NAND2X1 _12029_ (
    .A(_05580_),
    .B(_05581_),
    .Y(_05582_)
  );
  OAI22X1 _12030_ (
    .A(_05475_),
    .B(_05532_),
    .C(_05534_),
    .D(_05466_),
    .Y(_05583_)
  );
  NAND3X1 _12031_ (
    .A(_05580_),
    .B(_05581_),
    .C(_05583_),
    .Y(_05584_)
  );
  XOR2X1 _12032_ (
    .A(_05582_),
    .B(_05583_),
    .Y(_05585_)
  );
  XOR2X1 _12033_ (
    .A(_05574_),
    .B(_05585_),
    .Y(_05586_)
  );
  OAI21X1 _12034_ (
    .A(_05537_),
    .B(_05542_),
    .C(_05544_),
    .Y(_05587_)
  );
  NAND2X1 _12035_ (
    .A(multiplier_0.op1_7_ ),
    .B(_05276_),
    .Y(_05588_)
  );
  NOR2X1 _12036_ (
    .A(_05130_),
    .B(_05336_),
    .Y(_05589_)
  );
  NAND3X1 _12037_ (
    .A(multiplier_0.op1_5_ ),
    .B(_05303_),
    .C(_05589_),
    .Y(_05590_)
  );
  OAI21X1 _12038_ (
    .A(_05130_),
    .B(_05302_),
    .C(_05532_),
    .Y(_05591_)
  );
  NAND2X1 _12039_ (
    .A(_05590_),
    .B(_05591_),
    .Y(_05592_)
  );
  XOR2X1 _12040_ (
    .A(_05588_),
    .B(_05592_),
    .Y(_05593_)
  );
  AOI21X1 _12041_ (
    .A(_05538_),
    .B(_05539_),
    .C(_05541_),
    .Y(_05594_)
  );
  NAND2X1 _12042_ (
    .A(multiplier_0.op1_4_ ),
    .B(_05384_),
    .Y(_05595_)
  );
  NOR2X1 _12043_ (
    .A(_05127_),
    .B(_05429_),
    .Y(_05596_)
  );
  NOR2X1 _12044_ (
    .A(multiplier_0.op1_2_ ),
    .B(_05481_),
    .Y(_05597_)
  );
  AND2X1 _12045_ (
    .A(_05596_),
    .B(_05597_),
    .Y(_05598_)
  );
  XNOR2X1 _12046_ (
    .A(_05596_),
    .B(_05597_),
    .Y(_05599_)
  );
  NOR2X1 _12047_ (
    .A(_05595_),
    .B(_05599_),
    .Y(_05600_)
  );
  XNOR2X1 _12048_ (
    .A(_05595_),
    .B(_05599_),
    .Y(_05601_)
  );
  NOR2X1 _12049_ (
    .A(_05594_),
    .B(_05601_),
    .Y(_05602_)
  );
  XOR2X1 _12050_ (
    .A(_05594_),
    .B(_05601_),
    .Y(_05603_)
  );
  XOR2X1 _12051_ (
    .A(_05593_),
    .B(_05603_),
    .Y(_05604_)
  );
  AND2X1 _12052_ (
    .A(_05587_),
    .B(_05604_),
    .Y(_05605_)
  );
  XOR2X1 _12053_ (
    .A(_05587_),
    .B(_05604_),
    .Y(_05606_)
  );
  AND2X1 _12054_ (
    .A(_05586_),
    .B(_05606_),
    .Y(_05607_)
  );
  XNOR2X1 _12055_ (
    .A(_05586_),
    .B(_05606_),
    .Y(_05608_)
  );
  NOR2X1 _12056_ (
    .A(_05573_),
    .B(_05608_),
    .Y(_05609_)
  );
  XNOR2X1 _12057_ (
    .A(_05573_),
    .B(_05608_),
    .Y(_05610_)
  );
  AOI21X1 _12058_ (
    .A(_05526_),
    .B(_05529_),
    .C(_05610_),
    .Y(_05611_)
  );
  XNOR2X1 _12059_ (
    .A(_05571_),
    .B(_05610_),
    .Y(_05612_)
  );
  NAND2X1 _12060_ (
    .A(_05570_),
    .B(_05612_),
    .Y(_05613_)
  );
  XNOR2X1 _12061_ (
    .A(_05570_),
    .B(_05612_),
    .Y(_05614_)
  );
  NOR2X1 _12062_ (
    .A(_05553_),
    .B(_05614_),
    .Y(_05615_)
  );
  XOR2X1 _12063_ (
    .A(_05553_),
    .B(_05614_),
    .Y(_05616_)
  );
  OAI21X1 _12064_ (
    .A(_05511_),
    .B(_05558_),
    .C(_05556_),
    .Y(_05617_)
  );
  XNOR2X1 _12065_ (
    .A(_05616_),
    .B(_05617_),
    .Y(_05618_)
  );
  MUX2X1 _12066_ (
    .A(_05253_),
    .B(_05618_),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05619_)
  );
  NAND2X1 _12067_ (
    .A(multiplier_0.reslo_10_ ),
    .B(_05619_),
    .Y(_05620_)
  );
  XNOR2X1 _12068_ (
    .A(multiplier_0.reslo_10_ ),
    .B(_05619_),
    .Y(_05621_)
  );
  XNOR2X1 _12069_ (
    .A(_05569_),
    .B(_05621_),
    .Y(_05622_)
  );
  AND2X1 _12070_ (
    .A(_05225_),
    .B(_05622_),
    .Y(_05623_)
  );
  OAI21X1 _12071_ (
    .A(multiplier_0.reslo_10_ ),
    .B(_05225_),
    .C(_05222_),
    .Y(_05624_)
  );
  OR2X1 _12072_ (
    .A(_05183_),
    .B(_05219_),
    .Y(_05625_)
  );
  OAI21X1 _12073_ (
    .A(_05623_),
    .B(_05624_),
    .C(_05625_),
    .Y(_04448_)
  );
  OAI21X1 _12074_ (
    .A(_05569_),
    .B(_05621_),
    .C(_05620_),
    .Y(_05626_)
  );
  NOR2X1 _12075_ (
    .A(_05609_),
    .B(_05611_),
    .Y(_05627_)
  );
  OAI21X1 _12076_ (
    .A(_05574_),
    .B(_05585_),
    .C(_05584_),
    .Y(_05628_)
  );
  NOR2X1 _12077_ (
    .A(_05605_),
    .B(_05607_),
    .Y(_05629_)
  );
  OAI21X1 _12078_ (
    .A(_05575_),
    .B(_05579_),
    .C(_05578_),
    .Y(_05630_)
  );
  NAND2X1 _12079_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05212_),
    .Y(_05631_)
  );
  NAND2X1 _12080_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05230_),
    .Y(_05632_)
  );
  AND2X1 _12081_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05246_),
    .Y(_05633_)
  );
  NAND3X1 _12082_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05230_),
    .C(_05577_),
    .Y(_05634_)
  );
  XOR2X1 _12083_ (
    .A(_05577_),
    .B(_05632_),
    .Y(_05635_)
  );
  XNOR2X1 _12084_ (
    .A(_05631_),
    .B(_05635_),
    .Y(_05636_)
  );
  OAI21X1 _12085_ (
    .A(_05588_),
    .B(_05592_),
    .C(_05590_),
    .Y(_05637_)
  );
  INVX1 _12086_ (
    .A(_05637_),
    .Y(_05638_)
  );
  NOR2X1 _12087_ (
    .A(_05636_),
    .B(_05638_),
    .Y(_05639_)
  );
  XOR2X1 _12088_ (
    .A(_05636_),
    .B(_05637_),
    .Y(_05640_)
  );
  AOI21X1 _12089_ (
    .A(_05578_),
    .B(_05580_),
    .C(_05640_),
    .Y(_05641_)
  );
  XOR2X1 _12090_ (
    .A(_05630_),
    .B(_05640_),
    .Y(_05642_)
  );
  AOI21X1 _12091_ (
    .A(_05593_),
    .B(_05603_),
    .C(_05602_),
    .Y(_05643_)
  );
  NAND2X1 _12092_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05276_),
    .Y(_05644_)
  );
  NOR2X1 _12093_ (
    .A(_05131_),
    .B(_05302_),
    .Y(_05645_)
  );
  NAND2X1 _12094_ (
    .A(_05589_),
    .B(_05645_),
    .Y(_05646_)
  );
  XNOR2X1 _12095_ (
    .A(_05589_),
    .B(_05645_),
    .Y(_05647_)
  );
  XOR2X1 _12096_ (
    .A(_05644_),
    .B(_05647_),
    .Y(_05648_)
  );
  NOR2X1 _12097_ (
    .A(_05598_),
    .B(_05600_),
    .Y(_05649_)
  );
  NAND2X1 _12098_ (
    .A(multiplier_0.op1_5_ ),
    .B(_05384_),
    .Y(_05650_)
  );
  NOR2X1 _12099_ (
    .A(_05128_),
    .B(_05429_),
    .Y(_05651_)
  );
  NOR2X1 _12100_ (
    .A(multiplier_0.op1_3_ ),
    .B(_05481_),
    .Y(_05652_)
  );
  AND2X1 _12101_ (
    .A(_05651_),
    .B(_05652_),
    .Y(_05653_)
  );
  XNOR2X1 _12102_ (
    .A(_05651_),
    .B(_05652_),
    .Y(_05654_)
  );
  NOR2X1 _12103_ (
    .A(_05650_),
    .B(_05654_),
    .Y(_05655_)
  );
  XNOR2X1 _12104_ (
    .A(_05650_),
    .B(_05654_),
    .Y(_05656_)
  );
  INVX1 _12105_ (
    .A(_05656_),
    .Y(_05657_)
  );
  OAI21X1 _12106_ (
    .A(_05598_),
    .B(_05600_),
    .C(_05657_),
    .Y(_05658_)
  );
  XNOR2X1 _12107_ (
    .A(_05649_),
    .B(_05657_),
    .Y(_05659_)
  );
  NAND2X1 _12108_ (
    .A(_05648_),
    .B(_05659_),
    .Y(_05660_)
  );
  XOR2X1 _12109_ (
    .A(_05648_),
    .B(_05659_),
    .Y(_05661_)
  );
  INVX1 _12110_ (
    .A(_05661_),
    .Y(_05662_)
  );
  NOR2X1 _12111_ (
    .A(_05643_),
    .B(_05662_),
    .Y(_05663_)
  );
  XNOR2X1 _12112_ (
    .A(_05643_),
    .B(_05662_),
    .Y(_05664_)
  );
  NOR2X1 _12113_ (
    .A(_05642_),
    .B(_05664_),
    .Y(_05665_)
  );
  XOR2X1 _12114_ (
    .A(_05642_),
    .B(_05664_),
    .Y(_05666_)
  );
  OAI21X1 _12115_ (
    .A(_05605_),
    .B(_05607_),
    .C(_05666_),
    .Y(_05667_)
  );
  INVX1 _12116_ (
    .A(_05667_),
    .Y(_05668_)
  );
  XNOR2X1 _12117_ (
    .A(_05629_),
    .B(_05666_),
    .Y(_05669_)
  );
  XOR2X1 _12118_ (
    .A(_05628_),
    .B(_05669_),
    .Y(_05670_)
  );
  OAI21X1 _12119_ (
    .A(_05609_),
    .B(_05611_),
    .C(_05670_),
    .Y(_05671_)
  );
  XOR2X1 _12120_ (
    .A(_05627_),
    .B(_05670_),
    .Y(_05672_)
  );
  OR2X1 _12121_ (
    .A(_05613_),
    .B(_05672_),
    .Y(_05673_)
  );
  XNOR2X1 _12122_ (
    .A(_05613_),
    .B(_05672_),
    .Y(_05674_)
  );
  AOI21X1 _12123_ (
    .A(_05616_),
    .B(_05617_),
    .C(_05615_),
    .Y(_05675_)
  );
  XNOR2X1 _12124_ (
    .A(_05674_),
    .B(_05675_),
    .Y(_05676_)
  );
  MUX2X1 _12125_ (
    .A(_05281_),
    .B(_05676_),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05677_)
  );
  AND2X1 _12126_ (
    .A(multiplier_0.reslo_11_ ),
    .B(_05677_),
    .Y(_05678_)
  );
  XOR2X1 _12127_ (
    .A(multiplier_0.reslo_11_ ),
    .B(_05677_),
    .Y(_05679_)
  );
  XNOR2X1 _12128_ (
    .A(_05626_),
    .B(_05679_),
    .Y(_05680_)
  );
  OAI21X1 _12129_ (
    .A(multiplier_0.reslo_11_ ),
    .B(_05225_),
    .C(_05222_),
    .Y(_05681_)
  );
  AOI21X1 _12130_ (
    .A(_05225_),
    .B(_05680_),
    .C(_05681_),
    .Y(_05682_)
  );
  INVX1 _12131_ (
    .A(_05682_),
    .Y(_05683_)
  );
  OAI21X1 _12132_ (
    .A(_05185_),
    .B(_05219_),
    .C(_05683_),
    .Y(_04449_)
  );
  AOI21X1 _12133_ (
    .A(_05626_),
    .B(_05679_),
    .C(_05678_),
    .Y(_05684_)
  );
  OAI21X1 _12134_ (
    .A(_05674_),
    .B(_05675_),
    .C(_05673_),
    .Y(_05685_)
  );
  AOI21X1 _12135_ (
    .A(_05628_),
    .B(_05669_),
    .C(_05668_),
    .Y(_05686_)
  );
  NOR2X1 _12136_ (
    .A(_05639_),
    .B(_05641_),
    .Y(_05687_)
  );
  NOR2X1 _12137_ (
    .A(_05663_),
    .B(_05665_),
    .Y(_05688_)
  );
  OAI21X1 _12138_ (
    .A(_05631_),
    .B(_05635_),
    .C(_05634_),
    .Y(_05689_)
  );
  INVX1 _12139_ (
    .A(_05689_),
    .Y(_05690_)
  );
  NAND2X1 _12140_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05212_),
    .Y(_05691_)
  );
  NAND2X1 _12141_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05230_),
    .Y(_05692_)
  );
  AND2X1 _12142_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05246_),
    .Y(_05693_)
  );
  NAND3X1 _12143_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05230_),
    .C(_05633_),
    .Y(_05694_)
  );
  XOR2X1 _12144_ (
    .A(_05633_),
    .B(_05692_),
    .Y(_05695_)
  );
  XNOR2X1 _12145_ (
    .A(_05691_),
    .B(_05695_),
    .Y(_05696_)
  );
  OAI21X1 _12146_ (
    .A(_05644_),
    .B(_05647_),
    .C(_05646_),
    .Y(_05697_)
  );
  INVX1 _12147_ (
    .A(_05697_),
    .Y(_05698_)
  );
  NOR2X1 _12148_ (
    .A(_05696_),
    .B(_05698_),
    .Y(_05699_)
  );
  XOR2X1 _12149_ (
    .A(_05696_),
    .B(_05697_),
    .Y(_05700_)
  );
  NOR2X1 _12150_ (
    .A(_05690_),
    .B(_05700_),
    .Y(_05701_)
  );
  XNOR2X1 _12151_ (
    .A(_05689_),
    .B(_05700_),
    .Y(_05702_)
  );
  OAI21X1 _12152_ (
    .A(_05649_),
    .B(_05656_),
    .C(_05660_),
    .Y(_05703_)
  );
  NAND2X1 _12153_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05276_),
    .Y(_05704_)
  );
  NOR2X1 _12154_ (
    .A(_05132_),
    .B(_05336_),
    .Y(_05705_)
  );
  NAND2X1 _12155_ (
    .A(_05645_),
    .B(_05705_),
    .Y(_05706_)
  );
  OAI22X1 _12156_ (
    .A(_05132_),
    .B(_05302_),
    .C(_05336_),
    .D(_05131_),
    .Y(_05707_)
  );
  NAND2X1 _12157_ (
    .A(_05706_),
    .B(_05707_),
    .Y(_05708_)
  );
  XOR2X1 _12158_ (
    .A(_05704_),
    .B(_05708_),
    .Y(_05709_)
  );
  NOR2X1 _12159_ (
    .A(_05653_),
    .B(_05655_),
    .Y(_05710_)
  );
  NAND2X1 _12160_ (
    .A(multiplier_0.op1_6_ ),
    .B(_05384_),
    .Y(_05711_)
  );
  NOR2X1 _12161_ (
    .A(_05129_),
    .B(_05429_),
    .Y(_05712_)
  );
  NOR2X1 _12162_ (
    .A(multiplier_0.op1_4_ ),
    .B(_05481_),
    .Y(_05713_)
  );
  AND2X1 _12163_ (
    .A(_05712_),
    .B(_05713_),
    .Y(_05714_)
  );
  XNOR2X1 _12164_ (
    .A(_05712_),
    .B(_05713_),
    .Y(_05715_)
  );
  NOR2X1 _12165_ (
    .A(_05711_),
    .B(_05715_),
    .Y(_05716_)
  );
  XNOR2X1 _12166_ (
    .A(_05711_),
    .B(_05715_),
    .Y(_05717_)
  );
  INVX1 _12167_ (
    .A(_05717_),
    .Y(_05718_)
  );
  OAI21X1 _12168_ (
    .A(_05653_),
    .B(_05655_),
    .C(_05718_),
    .Y(_05719_)
  );
  XNOR2X1 _12169_ (
    .A(_05710_),
    .B(_05718_),
    .Y(_05720_)
  );
  NAND2X1 _12170_ (
    .A(_05709_),
    .B(_05720_),
    .Y(_05721_)
  );
  XNOR2X1 _12171_ (
    .A(_05709_),
    .B(_05720_),
    .Y(_05722_)
  );
  AOI21X1 _12172_ (
    .A(_05658_),
    .B(_05660_),
    .C(_05722_),
    .Y(_05723_)
  );
  XNOR2X1 _12173_ (
    .A(_05703_),
    .B(_05722_),
    .Y(_05724_)
  );
  AND2X1 _12174_ (
    .A(_05702_),
    .B(_05724_),
    .Y(_05725_)
  );
  NOR2X1 _12175_ (
    .A(_05702_),
    .B(_05724_),
    .Y(_05726_)
  );
  NOR2X1 _12176_ (
    .A(_05725_),
    .B(_05726_),
    .Y(_05727_)
  );
  OAI21X1 _12177_ (
    .A(_05663_),
    .B(_05665_),
    .C(_05727_),
    .Y(_05728_)
  );
  XNOR2X1 _12178_ (
    .A(_05688_),
    .B(_05727_),
    .Y(_05729_)
  );
  OAI21X1 _12179_ (
    .A(_05639_),
    .B(_05641_),
    .C(_05729_),
    .Y(_05730_)
  );
  XOR2X1 _12180_ (
    .A(_05687_),
    .B(_05729_),
    .Y(_05731_)
  );
  NOR2X1 _12181_ (
    .A(_05686_),
    .B(_05731_),
    .Y(_05732_)
  );
  XNOR2X1 _12182_ (
    .A(_05686_),
    .B(_05731_),
    .Y(_05733_)
  );
  NOR2X1 _12183_ (
    .A(_05671_),
    .B(_05733_),
    .Y(_05734_)
  );
  XOR2X1 _12184_ (
    .A(_05671_),
    .B(_05733_),
    .Y(_05735_)
  );
  XNOR2X1 _12185_ (
    .A(_05685_),
    .B(_05735_),
    .Y(_05736_)
  );
  NAND2X1 _12186_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05314_),
    .Y(_05737_)
  );
  OAI21X1 _12187_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05736_),
    .C(_05737_),
    .Y(_05738_)
  );
  NAND2X1 _12188_ (
    .A(multiplier_0.reslo_12_ ),
    .B(_05738_),
    .Y(_05739_)
  );
  XNOR2X1 _12189_ (
    .A(multiplier_0.reslo_12_ ),
    .B(_05738_),
    .Y(_05740_)
  );
  XOR2X1 _12190_ (
    .A(_05684_),
    .B(_05740_),
    .Y(_05741_)
  );
  NOR2X1 _12191_ (
    .A(multiplier_0.reslo_12_ ),
    .B(_05225_),
    .Y(_05742_)
  );
  NOR2X1 _12192_ (
    .A(_05221_),
    .B(_05742_),
    .Y(_05743_)
  );
  OAI21X1 _12193_ (
    .A(_05224_),
    .B(_05741_),
    .C(_05743_),
    .Y(_05744_)
  );
  OAI21X1 _12194_ (
    .A(_05187_),
    .B(_05219_),
    .C(_05744_),
    .Y(_04450_)
  );
  OAI21X1 _12195_ (
    .A(_05684_),
    .B(_05740_),
    .C(_05739_),
    .Y(_05745_)
  );
  AOI21X1 _12196_ (
    .A(_05685_),
    .B(_05735_),
    .C(_05734_),
    .Y(_05746_)
  );
  NAND2X1 _12197_ (
    .A(_05728_),
    .B(_05730_),
    .Y(_05747_)
  );
  NOR2X1 _12198_ (
    .A(_05699_),
    .B(_05701_),
    .Y(_05748_)
  );
  NOR2X1 _12199_ (
    .A(_05723_),
    .B(_05725_),
    .Y(_05749_)
  );
  OAI21X1 _12200_ (
    .A(_05691_),
    .B(_05695_),
    .C(_05694_),
    .Y(_05750_)
  );
  INVX1 _12201_ (
    .A(_05750_),
    .Y(_05751_)
  );
  NAND2X1 _12202_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05212_),
    .Y(_05752_)
  );
  NAND2X1 _12203_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05230_),
    .Y(_05753_)
  );
  AND2X1 _12204_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05246_),
    .Y(_05754_)
  );
  NAND3X1 _12205_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05230_),
    .C(_05693_),
    .Y(_05755_)
  );
  XOR2X1 _12206_ (
    .A(_05693_),
    .B(_05753_),
    .Y(_05756_)
  );
  XNOR2X1 _12207_ (
    .A(_05752_),
    .B(_05756_),
    .Y(_05757_)
  );
  OAI21X1 _12208_ (
    .A(_05704_),
    .B(_05708_),
    .C(_05706_),
    .Y(_05758_)
  );
  INVX1 _12209_ (
    .A(_05758_),
    .Y(_05759_)
  );
  NOR2X1 _12210_ (
    .A(_05757_),
    .B(_05759_),
    .Y(_05760_)
  );
  XOR2X1 _12211_ (
    .A(_05757_),
    .B(_05758_),
    .Y(_05761_)
  );
  NOR2X1 _12212_ (
    .A(_05751_),
    .B(_05761_),
    .Y(_05762_)
  );
  XNOR2X1 _12213_ (
    .A(_05750_),
    .B(_05761_),
    .Y(_05763_)
  );
  OAI21X1 _12214_ (
    .A(_05710_),
    .B(_05717_),
    .C(_05721_),
    .Y(_05764_)
  );
  NAND2X1 _12215_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05276_),
    .Y(_05765_)
  );
  AND2X1 _12216_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05303_),
    .Y(_05766_)
  );
  NAND2X1 _12217_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05337_),
    .Y(_05767_)
  );
  NAND2X1 _12218_ (
    .A(_05705_),
    .B(_05766_),
    .Y(_05768_)
  );
  XNOR2X1 _12219_ (
    .A(_05705_),
    .B(_05766_),
    .Y(_05769_)
  );
  XOR2X1 _12220_ (
    .A(_05765_),
    .B(_05769_),
    .Y(_05770_)
  );
  NOR2X1 _12221_ (
    .A(_05714_),
    .B(_05716_),
    .Y(_05771_)
  );
  NAND2X1 _12222_ (
    .A(multiplier_0.op1_7_ ),
    .B(_05384_),
    .Y(_05772_)
  );
  NOR2X1 _12223_ (
    .A(_05130_),
    .B(_05429_),
    .Y(_05773_)
  );
  NOR2X1 _12224_ (
    .A(multiplier_0.op1_5_ ),
    .B(_05481_),
    .Y(_05774_)
  );
  XNOR2X1 _12225_ (
    .A(_05773_),
    .B(_05774_),
    .Y(_05775_)
  );
  NOR2X1 _12226_ (
    .A(_05772_),
    .B(_05775_),
    .Y(_05776_)
  );
  XNOR2X1 _12227_ (
    .A(_05772_),
    .B(_05775_),
    .Y(_05777_)
  );
  INVX1 _12228_ (
    .A(_05777_),
    .Y(_05778_)
  );
  OAI21X1 _12229_ (
    .A(_05714_),
    .B(_05716_),
    .C(_05778_),
    .Y(_05779_)
  );
  XNOR2X1 _12230_ (
    .A(_05771_),
    .B(_05778_),
    .Y(_05780_)
  );
  NAND2X1 _12231_ (
    .A(_05770_),
    .B(_05780_),
    .Y(_05781_)
  );
  XNOR2X1 _12232_ (
    .A(_05770_),
    .B(_05780_),
    .Y(_05782_)
  );
  AOI21X1 _12233_ (
    .A(_05719_),
    .B(_05721_),
    .C(_05782_),
    .Y(_05783_)
  );
  XNOR2X1 _12234_ (
    .A(_05764_),
    .B(_05782_),
    .Y(_05784_)
  );
  AND2X1 _12235_ (
    .A(_05763_),
    .B(_05784_),
    .Y(_05785_)
  );
  NOR2X1 _12236_ (
    .A(_05763_),
    .B(_05784_),
    .Y(_05786_)
  );
  NOR2X1 _12237_ (
    .A(_05785_),
    .B(_05786_),
    .Y(_05787_)
  );
  OAI21X1 _12238_ (
    .A(_05723_),
    .B(_05725_),
    .C(_05787_),
    .Y(_05788_)
  );
  XNOR2X1 _12239_ (
    .A(_05749_),
    .B(_05787_),
    .Y(_05789_)
  );
  OAI21X1 _12240_ (
    .A(_05699_),
    .B(_05701_),
    .C(_05789_),
    .Y(_05790_)
  );
  XOR2X1 _12241_ (
    .A(_05748_),
    .B(_05789_),
    .Y(_05791_)
  );
  AOI21X1 _12242_ (
    .A(_05728_),
    .B(_05730_),
    .C(_05791_),
    .Y(_05792_)
  );
  XNOR2X1 _12243_ (
    .A(_05747_),
    .B(_05791_),
    .Y(_05793_)
  );
  NAND2X1 _12244_ (
    .A(_05732_),
    .B(_05793_),
    .Y(_05794_)
  );
  XNOR2X1 _12245_ (
    .A(_05732_),
    .B(_05793_),
    .Y(_05795_)
  );
  XOR2X1 _12246_ (
    .A(_05746_),
    .B(_05795_),
    .Y(_05796_)
  );
  NAND2X1 _12247_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05353_),
    .Y(_05797_)
  );
  OAI21X1 _12248_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05796_),
    .C(_05797_),
    .Y(_05798_)
  );
  NOR2X1 _12249_ (
    .A(_05138_),
    .B(_05798_),
    .Y(_05799_)
  );
  XNOR2X1 _12250_ (
    .A(multiplier_0.reslo_13_ ),
    .B(_05798_),
    .Y(_05800_)
  );
  XNOR2X1 _12251_ (
    .A(_05745_),
    .B(_05800_),
    .Y(_05801_)
  );
  OAI21X1 _12252_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.cycle_1_ ),
    .C(_05801_),
    .Y(_05802_)
  );
  NAND2X1 _12253_ (
    .A(_05138_),
    .B(_05224_),
    .Y(_05803_)
  );
  NAND3X1 _12254_ (
    .A(_05222_),
    .B(_05802_),
    .C(_05803_),
    .Y(_05804_)
  );
  OAI21X1 _12255_ (
    .A(_05189_),
    .B(_05219_),
    .C(_05804_),
    .Y(_04451_)
  );
  AOI21X1 _12256_ (
    .A(_05745_),
    .B(_05800_),
    .C(_05799_),
    .Y(_05805_)
  );
  OAI21X1 _12257_ (
    .A(_05746_),
    .B(_05795_),
    .C(_05794_),
    .Y(_05806_)
  );
  NAND2X1 _12258_ (
    .A(_05788_),
    .B(_05790_),
    .Y(_05807_)
  );
  NOR2X1 _12259_ (
    .A(_05760_),
    .B(_05762_),
    .Y(_05808_)
  );
  NOR2X1 _12260_ (
    .A(_05783_),
    .B(_05785_),
    .Y(_05809_)
  );
  OAI21X1 _12261_ (
    .A(_05752_),
    .B(_05756_),
    .C(_05755_),
    .Y(_05810_)
  );
  INVX1 _12262_ (
    .A(_05810_),
    .Y(_05811_)
  );
  NAND2X1 _12263_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05212_),
    .Y(_05812_)
  );
  NAND2X1 _12264_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05230_),
    .Y(_05813_)
  );
  AND2X1 _12265_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05246_),
    .Y(_05814_)
  );
  NAND3X1 _12266_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05230_),
    .C(_05754_),
    .Y(_05815_)
  );
  XOR2X1 _12267_ (
    .A(_05754_),
    .B(_05813_),
    .Y(_05816_)
  );
  XNOR2X1 _12268_ (
    .A(_05812_),
    .B(_05816_),
    .Y(_05817_)
  );
  OAI21X1 _12269_ (
    .A(_05765_),
    .B(_05769_),
    .C(_05768_),
    .Y(_05818_)
  );
  INVX1 _12270_ (
    .A(_05818_),
    .Y(_05819_)
  );
  NOR2X1 _12271_ (
    .A(_05817_),
    .B(_05819_),
    .Y(_05820_)
  );
  XOR2X1 _12272_ (
    .A(_05817_),
    .B(_05818_),
    .Y(_05821_)
  );
  NOR2X1 _12273_ (
    .A(_05811_),
    .B(_05821_),
    .Y(_05822_)
  );
  XNOR2X1 _12274_ (
    .A(_05810_),
    .B(_05821_),
    .Y(_05823_)
  );
  OAI21X1 _12275_ (
    .A(_05771_),
    .B(_05777_),
    .C(_05781_),
    .Y(_05824_)
  );
  NAND2X1 _12276_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05276_),
    .Y(_05825_)
  );
  AND2X1 _12277_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05303_),
    .Y(_05826_)
  );
  NAND2X1 _12278_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05337_),
    .Y(_05827_)
  );
  NAND3X1 _12279_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05337_),
    .C(_05826_),
    .Y(_05828_)
  );
  XOR2X1 _12280_ (
    .A(_05767_),
    .B(_05826_),
    .Y(_05829_)
  );
  XOR2X1 _12281_ (
    .A(_05825_),
    .B(_05829_),
    .Y(_05830_)
  );
  AOI21X1 _12282_ (
    .A(_05773_),
    .B(_05774_),
    .C(_05776_),
    .Y(_05831_)
  );
  NAND2X1 _12283_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05384_),
    .Y(_05832_)
  );
  NOR2X1 _12284_ (
    .A(_05131_),
    .B(_05429_),
    .Y(_05833_)
  );
  NOR2X1 _12285_ (
    .A(multiplier_0.op1_6_ ),
    .B(_05481_),
    .Y(_05834_)
  );
  AND2X1 _12286_ (
    .A(_05833_),
    .B(_05834_),
    .Y(_05835_)
  );
  XNOR2X1 _12287_ (
    .A(_05833_),
    .B(_05834_),
    .Y(_05836_)
  );
  NOR2X1 _12288_ (
    .A(_05832_),
    .B(_05836_),
    .Y(_05837_)
  );
  XNOR2X1 _12289_ (
    .A(_05832_),
    .B(_05836_),
    .Y(_05838_)
  );
  OR2X1 _12290_ (
    .A(_05831_),
    .B(_05838_),
    .Y(_05839_)
  );
  XOR2X1 _12291_ (
    .A(_05831_),
    .B(_05838_),
    .Y(_05840_)
  );
  NAND2X1 _12292_ (
    .A(_05830_),
    .B(_05840_),
    .Y(_05841_)
  );
  XNOR2X1 _12293_ (
    .A(_05830_),
    .B(_05840_),
    .Y(_05842_)
  );
  AOI21X1 _12294_ (
    .A(_05779_),
    .B(_05781_),
    .C(_05842_),
    .Y(_05843_)
  );
  XNOR2X1 _12295_ (
    .A(_05824_),
    .B(_05842_),
    .Y(_05844_)
  );
  AND2X1 _12296_ (
    .A(_05823_),
    .B(_05844_),
    .Y(_05845_)
  );
  NOR2X1 _12297_ (
    .A(_05823_),
    .B(_05844_),
    .Y(_05846_)
  );
  NOR2X1 _12298_ (
    .A(_05845_),
    .B(_05846_),
    .Y(_05847_)
  );
  OAI21X1 _12299_ (
    .A(_05783_),
    .B(_05785_),
    .C(_05847_),
    .Y(_05848_)
  );
  XNOR2X1 _12300_ (
    .A(_05809_),
    .B(_05847_),
    .Y(_05849_)
  );
  OAI21X1 _12301_ (
    .A(_05760_),
    .B(_05762_),
    .C(_05849_),
    .Y(_05850_)
  );
  XOR2X1 _12302_ (
    .A(_05808_),
    .B(_05849_),
    .Y(_05851_)
  );
  AOI21X1 _12303_ (
    .A(_05788_),
    .B(_05790_),
    .C(_05851_),
    .Y(_05852_)
  );
  XNOR2X1 _12304_ (
    .A(_05807_),
    .B(_05851_),
    .Y(_05853_)
  );
  NOR2X1 _12305_ (
    .A(_05792_),
    .B(_05853_),
    .Y(_05854_)
  );
  AND2X1 _12306_ (
    .A(_05792_),
    .B(_05853_),
    .Y(_05855_)
  );
  NOR2X1 _12307_ (
    .A(_05854_),
    .B(_05855_),
    .Y(_05856_)
  );
  XNOR2X1 _12308_ (
    .A(_05806_),
    .B(_05856_),
    .Y(_05857_)
  );
  NAND2X1 _12309_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05396_),
    .Y(_05858_)
  );
  OAI21X1 _12310_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05857_),
    .C(_05858_),
    .Y(_05859_)
  );
  NAND2X1 _12311_ (
    .A(multiplier_0.reslo_14_ ),
    .B(_05859_),
    .Y(_05860_)
  );
  NOR2X1 _12312_ (
    .A(multiplier_0.reslo_14_ ),
    .B(_05859_),
    .Y(_05861_)
  );
  XOR2X1 _12313_ (
    .A(multiplier_0.reslo_14_ ),
    .B(_05859_),
    .Y(_05862_)
  );
  XNOR2X1 _12314_ (
    .A(_05805_),
    .B(_05862_),
    .Y(_05863_)
  );
  NOR2X1 _12315_ (
    .A(_05224_),
    .B(_05863_),
    .Y(_04467_)
  );
  OAI21X1 _12316_ (
    .A(multiplier_0.reslo_14_ ),
    .B(_05225_),
    .C(_05222_),
    .Y(_04468_)
  );
  OAI22X1 _12317_ (
    .A(_05191_),
    .B(_05219_),
    .C(_04467_),
    .D(_04468_),
    .Y(_04452_)
  );
  OAI21X1 _12318_ (
    .A(_05805_),
    .B(_05861_),
    .C(_05860_),
    .Y(_04469_)
  );
  AOI21X1 _12319_ (
    .A(_05806_),
    .B(_05856_),
    .C(_05855_),
    .Y(_04470_)
  );
  NAND2X1 _12320_ (
    .A(_05848_),
    .B(_05850_),
    .Y(_04471_)
  );
  NOR2X1 _12321_ (
    .A(_05820_),
    .B(_05822_),
    .Y(_04472_)
  );
  NOR2X1 _12322_ (
    .A(_05843_),
    .B(_05845_),
    .Y(_04473_)
  );
  OAI21X1 _12323_ (
    .A(_05812_),
    .B(_05816_),
    .C(_05815_),
    .Y(_04474_)
  );
  INVX1 _12324_ (
    .A(_04474_),
    .Y(_04475_)
  );
  NAND2X1 _12325_ (
    .A(multiplier_0.op1_15_ ),
    .B(_05212_),
    .Y(_04476_)
  );
  NAND2X1 _12326_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05230_),
    .Y(_04477_)
  );
  NAND3X1 _12327_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05230_),
    .C(_05814_),
    .Y(_04478_)
  );
  XOR2X1 _12328_ (
    .A(_05814_),
    .B(_04477_),
    .Y(_04479_)
  );
  XNOR2X1 _12329_ (
    .A(_04476_),
    .B(_04479_),
    .Y(_04480_)
  );
  OAI21X1 _12330_ (
    .A(_05825_),
    .B(_05829_),
    .C(_05828_),
    .Y(_04481_)
  );
  INVX1 _12331_ (
    .A(_04481_),
    .Y(_04482_)
  );
  NOR2X1 _12332_ (
    .A(_04480_),
    .B(_04482_),
    .Y(_04483_)
  );
  XOR2X1 _12333_ (
    .A(_04480_),
    .B(_04481_),
    .Y(_04484_)
  );
  NOR2X1 _12334_ (
    .A(_04475_),
    .B(_04484_),
    .Y(_04485_)
  );
  XNOR2X1 _12335_ (
    .A(_04474_),
    .B(_04484_),
    .Y(_04486_)
  );
  OAI21X1 _12336_ (
    .A(_05831_),
    .B(_05838_),
    .C(_05841_),
    .Y(_04487_)
  );
  NAND2X1 _12337_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05276_),
    .Y(_04488_)
  );
  AND2X1 _12338_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05303_),
    .Y(_04489_)
  );
  NAND2X1 _12339_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05337_),
    .Y(_04490_)
  );
  NAND3X1 _12340_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05337_),
    .C(_04489_),
    .Y(_04491_)
  );
  XOR2X1 _12341_ (
    .A(_05827_),
    .B(_04489_),
    .Y(_04492_)
  );
  XOR2X1 _12342_ (
    .A(_04488_),
    .B(_04492_),
    .Y(_04493_)
  );
  NOR2X1 _12343_ (
    .A(_05835_),
    .B(_05837_),
    .Y(_04494_)
  );
  NAND2X1 _12344_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05384_),
    .Y(_04495_)
  );
  NOR2X1 _12345_ (
    .A(_05132_),
    .B(_05429_),
    .Y(_04496_)
  );
  NOR2X1 _12346_ (
    .A(multiplier_0.op1_7_ ),
    .B(_05481_),
    .Y(_04497_)
  );
  XNOR2X1 _12347_ (
    .A(_04496_),
    .B(_04497_),
    .Y(_04498_)
  );
  NOR2X1 _12348_ (
    .A(_04495_),
    .B(_04498_),
    .Y(_04499_)
  );
  XNOR2X1 _12349_ (
    .A(_04495_),
    .B(_04498_),
    .Y(_04500_)
  );
  INVX1 _12350_ (
    .A(_04500_),
    .Y(_04501_)
  );
  OAI21X1 _12351_ (
    .A(_05835_),
    .B(_05837_),
    .C(_04501_),
    .Y(_04502_)
  );
  XNOR2X1 _12352_ (
    .A(_04494_),
    .B(_04501_),
    .Y(_04503_)
  );
  NAND2X1 _12353_ (
    .A(_04493_),
    .B(_04503_),
    .Y(_04504_)
  );
  XNOR2X1 _12354_ (
    .A(_04493_),
    .B(_04503_),
    .Y(_04505_)
  );
  AOI21X1 _12355_ (
    .A(_05839_),
    .B(_05841_),
    .C(_04505_),
    .Y(_04506_)
  );
  XNOR2X1 _12356_ (
    .A(_04487_),
    .B(_04505_),
    .Y(_04507_)
  );
  AND2X1 _12357_ (
    .A(_04486_),
    .B(_04507_),
    .Y(_04508_)
  );
  NOR2X1 _12358_ (
    .A(_04486_),
    .B(_04507_),
    .Y(_04509_)
  );
  NOR2X1 _12359_ (
    .A(_04508_),
    .B(_04509_),
    .Y(_04510_)
  );
  OAI21X1 _12360_ (
    .A(_05843_),
    .B(_05845_),
    .C(_04510_),
    .Y(_04511_)
  );
  XNOR2X1 _12361_ (
    .A(_04473_),
    .B(_04510_),
    .Y(_04512_)
  );
  OAI21X1 _12362_ (
    .A(_05820_),
    .B(_05822_),
    .C(_04512_),
    .Y(_04513_)
  );
  XOR2X1 _12363_ (
    .A(_04472_),
    .B(_04512_),
    .Y(_04514_)
  );
  AOI21X1 _12364_ (
    .A(_05848_),
    .B(_05850_),
    .C(_04514_),
    .Y(_04515_)
  );
  XNOR2X1 _12365_ (
    .A(_04471_),
    .B(_04514_),
    .Y(_04516_)
  );
  NAND2X1 _12366_ (
    .A(_05852_),
    .B(_04516_),
    .Y(_04517_)
  );
  XNOR2X1 _12367_ (
    .A(_05852_),
    .B(_04516_),
    .Y(_04518_)
  );
  XOR2X1 _12368_ (
    .A(_04470_),
    .B(_04518_),
    .Y(_04519_)
  );
  NAND2X1 _12369_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05448_),
    .Y(_04520_)
  );
  OAI21X1 _12370_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04519_),
    .C(_04520_),
    .Y(_04521_)
  );
  NOR2X1 _12371_ (
    .A(_05139_),
    .B(_04521_),
    .Y(_04522_)
  );
  XNOR2X1 _12372_ (
    .A(multiplier_0.reslo_15_ ),
    .B(_04521_),
    .Y(_04523_)
  );
  XNOR2X1 _12373_ (
    .A(_04469_),
    .B(_04523_),
    .Y(_04524_)
  );
  OAI21X1 _12374_ (
    .A(multiplier_0.reslo_15_ ),
    .B(_05225_),
    .C(_05222_),
    .Y(_04525_)
  );
  AOI21X1 _12375_ (
    .A(_05225_),
    .B(_04524_),
    .C(_04525_),
    .Y(_04526_)
  );
  INVX1 _12376_ (
    .A(_04526_),
    .Y(_04527_)
  );
  OAI21X1 _12377_ (
    .A(_05193_),
    .B(_05219_),
    .C(_04527_),
    .Y(_04453_)
  );
  AOI21X1 _12378_ (
    .A(_04469_),
    .B(_04523_),
    .C(_04522_),
    .Y(_04528_)
  );
  OAI21X1 _12379_ (
    .A(_04470_),
    .B(_04518_),
    .C(_04517_),
    .Y(_04529_)
  );
  NAND2X1 _12380_ (
    .A(_04511_),
    .B(_04513_),
    .Y(_04530_)
  );
  NOR2X1 _12381_ (
    .A(_04483_),
    .B(_04485_),
    .Y(_04531_)
  );
  NOR2X1 _12382_ (
    .A(_04506_),
    .B(_04508_),
    .Y(_04532_)
  );
  OAI21X1 _12383_ (
    .A(_04476_),
    .B(_04479_),
    .C(_04478_),
    .Y(_04533_)
  );
  INVX1 _12384_ (
    .A(_04533_),
    .Y(_04534_)
  );
  AND2X1 _12385_ (
    .A(multiplier_0.op1_15_ ),
    .B(multiplier_0.sign_sel ),
    .Y(_04535_)
  );
  NAND2X1 _12386_ (
    .A(multiplier_0.op1_15_ ),
    .B(multiplier_0.sign_sel ),
    .Y(_04536_)
  );
  NOR2X1 _12387_ (
    .A(_05213_),
    .B(_04536_),
    .Y(_04537_)
  );
  NAND2X1 _12388_ (
    .A(_05212_),
    .B(_04535_),
    .Y(_04538_)
  );
  NAND2X1 _12389_ (
    .A(multiplier_0.op1_15_ ),
    .B(_05230_),
    .Y(_04539_)
  );
  NAND2X1 _12390_ (
    .A(multiplier_0.op1_15_ ),
    .B(_05246_),
    .Y(_04540_)
  );
  OAI21X1 _12391_ (
    .A(_05133_),
    .B(_05245_),
    .C(_04539_),
    .Y(_04541_)
  );
  OAI21X1 _12392_ (
    .A(_04477_),
    .B(_04540_),
    .C(_04541_),
    .Y(_04542_)
  );
  XNOR2X1 _12393_ (
    .A(_04538_),
    .B(_04542_),
    .Y(_04543_)
  );
  OAI21X1 _12394_ (
    .A(_04488_),
    .B(_04492_),
    .C(_04491_),
    .Y(_04544_)
  );
  INVX1 _12395_ (
    .A(_04544_),
    .Y(_04545_)
  );
  NOR2X1 _12396_ (
    .A(_04543_),
    .B(_04545_),
    .Y(_04546_)
  );
  XNOR2X1 _12397_ (
    .A(_04543_),
    .B(_04545_),
    .Y(_04547_)
  );
  NOR2X1 _12398_ (
    .A(_04534_),
    .B(_04547_),
    .Y(_04548_)
  );
  XNOR2X1 _12399_ (
    .A(_04533_),
    .B(_04547_),
    .Y(_04549_)
  );
  OAI21X1 _12400_ (
    .A(_04494_),
    .B(_04500_),
    .C(_04504_),
    .Y(_04550_)
  );
  NAND2X1 _12401_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05276_),
    .Y(_04551_)
  );
  AND2X1 _12402_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05303_),
    .Y(_04552_)
  );
  NAND2X1 _12403_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05337_),
    .Y(_04553_)
  );
  NAND3X1 _12404_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05337_),
    .C(_04552_),
    .Y(_04554_)
  );
  XOR2X1 _12405_ (
    .A(_04490_),
    .B(_04552_),
    .Y(_04555_)
  );
  XOR2X1 _12406_ (
    .A(_04551_),
    .B(_04555_),
    .Y(_04556_)
  );
  AOI21X1 _12407_ (
    .A(_04496_),
    .B(_04497_),
    .C(_04499_),
    .Y(_04557_)
  );
  NAND2X1 _12408_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05384_),
    .Y(_04558_)
  );
  AND2X1 _12409_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05430_),
    .Y(_04559_)
  );
  NOR2X1 _12410_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05481_),
    .Y(_04560_)
  );
  XNOR2X1 _12411_ (
    .A(_04559_),
    .B(_04560_),
    .Y(_04561_)
  );
  NOR2X1 _12412_ (
    .A(_04558_),
    .B(_04561_),
    .Y(_04562_)
  );
  XNOR2X1 _12413_ (
    .A(_04558_),
    .B(_04561_),
    .Y(_04563_)
  );
  NOR2X1 _12414_ (
    .A(_04557_),
    .B(_04563_),
    .Y(_04564_)
  );
  XOR2X1 _12415_ (
    .A(_04557_),
    .B(_04563_),
    .Y(_04565_)
  );
  XNOR2X1 _12416_ (
    .A(_04556_),
    .B(_04565_),
    .Y(_04566_)
  );
  AOI21X1 _12417_ (
    .A(_04502_),
    .B(_04504_),
    .C(_04566_),
    .Y(_04567_)
  );
  XNOR2X1 _12418_ (
    .A(_04550_),
    .B(_04566_),
    .Y(_04568_)
  );
  AND2X1 _12419_ (
    .A(_04549_),
    .B(_04568_),
    .Y(_04569_)
  );
  NOR2X1 _12420_ (
    .A(_04549_),
    .B(_04568_),
    .Y(_04570_)
  );
  NOR2X1 _12421_ (
    .A(_04569_),
    .B(_04570_),
    .Y(_04571_)
  );
  OAI21X1 _12422_ (
    .A(_04506_),
    .B(_04508_),
    .C(_04571_),
    .Y(_04572_)
  );
  XNOR2X1 _12423_ (
    .A(_04532_),
    .B(_04571_),
    .Y(_04573_)
  );
  OAI21X1 _12424_ (
    .A(_04483_),
    .B(_04485_),
    .C(_04573_),
    .Y(_04574_)
  );
  XOR2X1 _12425_ (
    .A(_04531_),
    .B(_04573_),
    .Y(_04575_)
  );
  AOI21X1 _12426_ (
    .A(_04511_),
    .B(_04513_),
    .C(_04575_),
    .Y(_04576_)
  );
  XNOR2X1 _12427_ (
    .A(_04530_),
    .B(_04575_),
    .Y(_04577_)
  );
  AND2X1 _12428_ (
    .A(_04515_),
    .B(_04577_),
    .Y(_04578_)
  );
  NOR2X1 _12429_ (
    .A(_04515_),
    .B(_04577_),
    .Y(_04579_)
  );
  NOR2X1 _12430_ (
    .A(_04578_),
    .B(_04579_),
    .Y(_04580_)
  );
  XNOR2X1 _12431_ (
    .A(_04529_),
    .B(_04580_),
    .Y(_04581_)
  );
  MUX2X1 _12432_ (
    .A(_05503_),
    .B(_04581_),
    .S(multiplier_0.cycle_0_ ),
    .Y(_04582_)
  );
  NAND2X1 _12433_ (
    .A(multiplier_0.reshi_0_ ),
    .B(_04582_),
    .Y(_04583_)
  );
  NOR2X1 _12434_ (
    .A(multiplier_0.reshi_0_ ),
    .B(_04582_),
    .Y(_04584_)
  );
  XOR2X1 _12435_ (
    .A(multiplier_0.reshi_0_ ),
    .B(_04582_),
    .Y(_04585_)
  );
  XNOR2X1 _12436_ (
    .A(_04528_),
    .B(_04585_),
    .Y(_04586_)
  );
  NOR2X1 _12437_ (
    .A(multiplier_0.reshi_0_ ),
    .B(_05225_),
    .Y(_04587_)
  );
  NAND3X1 _12438_ (
    .A(_00101_),
    .B(_05103_),
    .C(_00102_),
    .Y(_04588_)
  );
  OR2X1 _12439_ (
    .A(_05168_),
    .B(_04588_),
    .Y(_04589_)
  );
  OAI21X1 _12440_ (
    .A(multiplier_0.acc_sel ),
    .B(_05169_),
    .C(_04589_),
    .Y(_04590_)
  );
  INVX1 _12441_ (
    .A(_04590_),
    .Y(_04591_)
  );
  OAI21X1 _12442_ (
    .A(_05224_),
    .B(_04586_),
    .C(_04591_),
    .Y(_04592_)
  );
  OAI22X1 _12443_ (
    .A(_05109_),
    .B(_04589_),
    .C(_04592_),
    .D(_04587_),
    .Y(_04431_)
  );
  OAI21X1 _12444_ (
    .A(_04528_),
    .B(_04584_),
    .C(_04583_),
    .Y(_04593_)
  );
  AOI21X1 _12445_ (
    .A(_04529_),
    .B(_04580_),
    .C(_04578_),
    .Y(_04594_)
  );
  NAND2X1 _12446_ (
    .A(_04572_),
    .B(_04574_),
    .Y(_04595_)
  );
  NOR2X1 _12447_ (
    .A(_04546_),
    .B(_04548_),
    .Y(_04596_)
  );
  NOR2X1 _12448_ (
    .A(_04567_),
    .B(_04569_),
    .Y(_04597_)
  );
  OAI22X1 _12449_ (
    .A(_04477_),
    .B(_04540_),
    .C(_04542_),
    .D(_04538_),
    .Y(_04598_)
  );
  OAI21X1 _12450_ (
    .A(_04551_),
    .B(_04555_),
    .C(_04554_),
    .Y(_04599_)
  );
  INVX1 _12451_ (
    .A(_04599_),
    .Y(_04600_)
  );
  NAND3X1 _12452_ (
    .A(_05230_),
    .B(_05246_),
    .C(_04535_),
    .Y(_04601_)
  );
  OAI21X1 _12453_ (
    .A(_05229_),
    .B(_04536_),
    .C(_04540_),
    .Y(_04602_)
  );
  NAND2X1 _12454_ (
    .A(_04601_),
    .B(_04602_),
    .Y(_04603_)
  );
  XNOR2X1 _12455_ (
    .A(_04538_),
    .B(_04603_),
    .Y(_04604_)
  );
  XNOR2X1 _12456_ (
    .A(_04599_),
    .B(_04604_),
    .Y(_04605_)
  );
  NAND2X1 _12457_ (
    .A(_04598_),
    .B(_04605_),
    .Y(_04606_)
  );
  XNOR2X1 _12458_ (
    .A(_04598_),
    .B(_04605_),
    .Y(_04607_)
  );
  INVX1 _12459_ (
    .A(_04607_),
    .Y(_04608_)
  );
  AOI21X1 _12460_ (
    .A(_04556_),
    .B(_04565_),
    .C(_04564_),
    .Y(_04609_)
  );
  NOR2X1 _12461_ (
    .A(_05133_),
    .B(_05275_),
    .Y(_04610_)
  );
  AND2X1 _12462_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05303_),
    .Y(_04611_)
  );
  NAND2X1 _12463_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05337_),
    .Y(_04612_)
  );
  NAND3X1 _12464_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05337_),
    .C(_04611_),
    .Y(_04613_)
  );
  XOR2X1 _12465_ (
    .A(_04553_),
    .B(_04611_),
    .Y(_04614_)
  );
  INVX1 _12466_ (
    .A(_04614_),
    .Y(_04615_)
  );
  NAND2X1 _12467_ (
    .A(_04610_),
    .B(_04615_),
    .Y(_04616_)
  );
  XNOR2X1 _12468_ (
    .A(_04610_),
    .B(_04614_),
    .Y(_04617_)
  );
  AOI21X1 _12469_ (
    .A(_04559_),
    .B(_04560_),
    .C(_04562_),
    .Y(_04618_)
  );
  NAND2X1 _12470_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05384_),
    .Y(_04619_)
  );
  AND2X1 _12471_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05430_),
    .Y(_04620_)
  );
  NOR2X1 _12472_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05481_),
    .Y(_04621_)
  );
  XNOR2X1 _12473_ (
    .A(_04620_),
    .B(_04621_),
    .Y(_04622_)
  );
  NOR2X1 _12474_ (
    .A(_04619_),
    .B(_04622_),
    .Y(_04623_)
  );
  XNOR2X1 _12475_ (
    .A(_04619_),
    .B(_04622_),
    .Y(_04624_)
  );
  NOR2X1 _12476_ (
    .A(_04618_),
    .B(_04624_),
    .Y(_04625_)
  );
  XOR2X1 _12477_ (
    .A(_04618_),
    .B(_04624_),
    .Y(_04626_)
  );
  XOR2X1 _12478_ (
    .A(_04617_),
    .B(_04626_),
    .Y(_04627_)
  );
  INVX1 _12479_ (
    .A(_04627_),
    .Y(_04628_)
  );
  NOR2X1 _12480_ (
    .A(_04609_),
    .B(_04628_),
    .Y(_04629_)
  );
  XNOR2X1 _12481_ (
    .A(_04609_),
    .B(_04627_),
    .Y(_04630_)
  );
  XNOR2X1 _12482_ (
    .A(_04607_),
    .B(_04630_),
    .Y(_04631_)
  );
  OAI21X1 _12483_ (
    .A(_04567_),
    .B(_04569_),
    .C(_04631_),
    .Y(_04632_)
  );
  XNOR2X1 _12484_ (
    .A(_04597_),
    .B(_04631_),
    .Y(_04633_)
  );
  OAI21X1 _12485_ (
    .A(_04546_),
    .B(_04548_),
    .C(_04633_),
    .Y(_04634_)
  );
  XOR2X1 _12486_ (
    .A(_04596_),
    .B(_04633_),
    .Y(_04635_)
  );
  AOI21X1 _12487_ (
    .A(_04572_),
    .B(_04574_),
    .C(_04635_),
    .Y(_04636_)
  );
  XNOR2X1 _12488_ (
    .A(_04595_),
    .B(_04635_),
    .Y(_04637_)
  );
  NAND2X1 _12489_ (
    .A(_04576_),
    .B(_04637_),
    .Y(_04638_)
  );
  XNOR2X1 _12490_ (
    .A(_04576_),
    .B(_04637_),
    .Y(_04639_)
  );
  XOR2X1 _12491_ (
    .A(_04594_),
    .B(_04639_),
    .Y(_04640_)
  );
  NAND2X1 _12492_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05560_),
    .Y(_04641_)
  );
  OAI21X1 _12493_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04640_),
    .C(_04641_),
    .Y(_04642_)
  );
  NAND2X1 _12494_ (
    .A(_05140_),
    .B(_04642_),
    .Y(_04643_)
  );
  NOR2X1 _12495_ (
    .A(_05140_),
    .B(_04642_),
    .Y(_04644_)
  );
  XNOR2X1 _12496_ (
    .A(multiplier_0.reshi_1_ ),
    .B(_04642_),
    .Y(_04645_)
  );
  XNOR2X1 _12497_ (
    .A(_04593_),
    .B(_04645_),
    .Y(_04646_)
  );
  AOI21X1 _12498_ (
    .A(_05225_),
    .B(_04646_),
    .C(_04590_),
    .Y(_04647_)
  );
  OAI21X1 _12499_ (
    .A(multiplier_0.reshi_1_ ),
    .B(_05225_),
    .C(_04647_),
    .Y(_04648_)
  );
  OAI21X1 _12500_ (
    .A(_05111_),
    .B(_04589_),
    .C(_04648_),
    .Y(_04438_)
  );
  OAI21X1 _12501_ (
    .A(_04594_),
    .B(_04639_),
    .C(_04638_),
    .Y(_04649_)
  );
  NAND2X1 _12502_ (
    .A(_04632_),
    .B(_04634_),
    .Y(_04650_)
  );
  OAI21X1 _12503_ (
    .A(_04600_),
    .B(_04604_),
    .C(_04606_),
    .Y(_04651_)
  );
  AOI21X1 _12504_ (
    .A(_04608_),
    .B(_04630_),
    .C(_04629_),
    .Y(_04652_)
  );
  INVX1 _12505_ (
    .A(_04652_),
    .Y(_04653_)
  );
  OAI21X1 _12506_ (
    .A(_04538_),
    .B(_04603_),
    .C(_04601_),
    .Y(_04654_)
  );
  NAND2X1 _12507_ (
    .A(_04613_),
    .B(_04616_),
    .Y(_04655_)
  );
  OAI21X1 _12508_ (
    .A(_05230_),
    .B(_05246_),
    .C(_04535_),
    .Y(_04656_)
  );
  NOR2X1 _12509_ (
    .A(_04654_),
    .B(_04656_),
    .Y(_04657_)
  );
  AOI21X1 _12510_ (
    .A(_04537_),
    .B(_04603_),
    .C(_04657_),
    .Y(_04658_)
  );
  AOI21X1 _12511_ (
    .A(_04613_),
    .B(_04616_),
    .C(_04658_),
    .Y(_04659_)
  );
  XNOR2X1 _12512_ (
    .A(_04655_),
    .B(_04658_),
    .Y(_04660_)
  );
  XOR2X1 _12513_ (
    .A(_04654_),
    .B(_04660_),
    .Y(_04661_)
  );
  AOI21X1 _12514_ (
    .A(_04617_),
    .B(_04626_),
    .C(_04625_),
    .Y(_04662_)
  );
  AND2X1 _12515_ (
    .A(multiplier_0.op1_15_ ),
    .B(_05276_),
    .Y(_04663_)
  );
  NAND2X1 _12516_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05303_),
    .Y(_04664_)
  );
  OR2X1 _12517_ (
    .A(_04612_),
    .B(_04664_),
    .Y(_04665_)
  );
  XNOR2X1 _12518_ (
    .A(_04612_),
    .B(_04664_),
    .Y(_04666_)
  );
  INVX1 _12519_ (
    .A(_04666_),
    .Y(_04667_)
  );
  NAND2X1 _12520_ (
    .A(_04663_),
    .B(_04667_),
    .Y(_04668_)
  );
  XNOR2X1 _12521_ (
    .A(_04663_),
    .B(_04666_),
    .Y(_04669_)
  );
  AOI21X1 _12522_ (
    .A(_04620_),
    .B(_04621_),
    .C(_04623_),
    .Y(_04670_)
  );
  NAND2X1 _12523_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05384_),
    .Y(_04671_)
  );
  AND2X1 _12524_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05430_),
    .Y(_04672_)
  );
  NOR2X1 _12525_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05481_),
    .Y(_04673_)
  );
  XNOR2X1 _12526_ (
    .A(_04672_),
    .B(_04673_),
    .Y(_04674_)
  );
  NOR2X1 _12527_ (
    .A(_04671_),
    .B(_04674_),
    .Y(_04675_)
  );
  XNOR2X1 _12528_ (
    .A(_04671_),
    .B(_04674_),
    .Y(_04676_)
  );
  NOR2X1 _12529_ (
    .A(_04670_),
    .B(_04676_),
    .Y(_04677_)
  );
  XOR2X1 _12530_ (
    .A(_04670_),
    .B(_04676_),
    .Y(_04678_)
  );
  XOR2X1 _12531_ (
    .A(_04669_),
    .B(_04678_),
    .Y(_04679_)
  );
  INVX1 _12532_ (
    .A(_04679_),
    .Y(_04680_)
  );
  NOR2X1 _12533_ (
    .A(_04662_),
    .B(_04680_),
    .Y(_04681_)
  );
  XNOR2X1 _12534_ (
    .A(_04662_),
    .B(_04679_),
    .Y(_04682_)
  );
  XOR2X1 _12535_ (
    .A(_04661_),
    .B(_04682_),
    .Y(_04683_)
  );
  NAND2X1 _12536_ (
    .A(_04653_),
    .B(_04683_),
    .Y(_04684_)
  );
  XNOR2X1 _12537_ (
    .A(_04652_),
    .B(_04683_),
    .Y(_04685_)
  );
  NAND2X1 _12538_ (
    .A(_04651_),
    .B(_04685_),
    .Y(_04686_)
  );
  XNOR2X1 _12539_ (
    .A(_04651_),
    .B(_04685_),
    .Y(_04687_)
  );
  AOI21X1 _12540_ (
    .A(_04632_),
    .B(_04634_),
    .C(_04687_),
    .Y(_04688_)
  );
  XNOR2X1 _12541_ (
    .A(_04650_),
    .B(_04687_),
    .Y(_04689_)
  );
  AND2X1 _12542_ (
    .A(_04636_),
    .B(_04689_),
    .Y(_04690_)
  );
  NOR2X1 _12543_ (
    .A(_04636_),
    .B(_04689_),
    .Y(_04691_)
  );
  NOR2X1 _12544_ (
    .A(_04690_),
    .B(_04691_),
    .Y(_04692_)
  );
  XNOR2X1 _12545_ (
    .A(_04649_),
    .B(_04692_),
    .Y(_04693_)
  );
  MUX2X1 _12546_ (
    .A(_05618_),
    .B(_04693_),
    .S(multiplier_0.cycle_0_ ),
    .Y(_04694_)
  );
  NAND2X1 _12547_ (
    .A(multiplier_0.reshi_2_ ),
    .B(_04694_),
    .Y(_04695_)
  );
  XNOR2X1 _12548_ (
    .A(multiplier_0.reshi_2_ ),
    .B(_04694_),
    .Y(_04696_)
  );
  AOI21X1 _12549_ (
    .A(_04593_),
    .B(_04643_),
    .C(_04644_),
    .Y(_04697_)
  );
  XNOR2X1 _12550_ (
    .A(_04696_),
    .B(_04697_),
    .Y(_04698_)
  );
  AOI21X1 _12551_ (
    .A(_05225_),
    .B(_04698_),
    .C(_04590_),
    .Y(_04699_)
  );
  OAI21X1 _12552_ (
    .A(multiplier_0.reshi_2_ ),
    .B(_05225_),
    .C(_04699_),
    .Y(_04700_)
  );
  OAI21X1 _12553_ (
    .A(_05113_),
    .B(_04589_),
    .C(_04700_),
    .Y(_04439_)
  );
  OAI21X1 _12554_ (
    .A(_04696_),
    .B(_04697_),
    .C(_04695_),
    .Y(_04701_)
  );
  AOI21X1 _12555_ (
    .A(_04649_),
    .B(_04692_),
    .C(_04690_),
    .Y(_04702_)
  );
  NAND2X1 _12556_ (
    .A(_04684_),
    .B(_04686_),
    .Y(_04703_)
  );
  AOI21X1 _12557_ (
    .A(_04654_),
    .B(_04660_),
    .C(_04659_),
    .Y(_04704_)
  );
  INVX1 _12558_ (
    .A(_04704_),
    .Y(_04705_)
  );
  AOI21X1 _12559_ (
    .A(_04661_),
    .B(_04682_),
    .C(_04681_),
    .Y(_04706_)
  );
  INVX1 _12560_ (
    .A(_04706_),
    .Y(_04707_)
  );
  OAI21X1 _12561_ (
    .A(_04612_),
    .B(_04664_),
    .C(_04668_),
    .Y(_04708_)
  );
  AOI21X1 _12562_ (
    .A(_04665_),
    .B(_04668_),
    .C(_04658_),
    .Y(_04709_)
  );
  XNOR2X1 _12563_ (
    .A(_04658_),
    .B(_04708_),
    .Y(_04710_)
  );
  XOR2X1 _12564_ (
    .A(_04654_),
    .B(_04710_),
    .Y(_04711_)
  );
  AOI21X1 _12565_ (
    .A(_04669_),
    .B(_04678_),
    .C(_04677_),
    .Y(_04712_)
  );
  NOR2X1 _12566_ (
    .A(_05275_),
    .B(_04536_),
    .Y(_04713_)
  );
  NAND2X1 _12567_ (
    .A(_05276_),
    .B(_04535_),
    .Y(_04714_)
  );
  NAND2X1 _12568_ (
    .A(multiplier_0.op1_15_ ),
    .B(_05303_),
    .Y(_04715_)
  );
  NAND2X1 _12569_ (
    .A(multiplier_0.op1_15_ ),
    .B(_05337_),
    .Y(_04716_)
  );
  OAI21X1 _12570_ (
    .A(_05133_),
    .B(_05336_),
    .C(_04715_),
    .Y(_04717_)
  );
  OAI21X1 _12571_ (
    .A(_04664_),
    .B(_04716_),
    .C(_04717_),
    .Y(_04718_)
  );
  XNOR2X1 _12572_ (
    .A(_04713_),
    .B(_04718_),
    .Y(_04719_)
  );
  AOI21X1 _12573_ (
    .A(_04672_),
    .B(_04673_),
    .C(_04675_),
    .Y(_04720_)
  );
  NAND2X1 _12574_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05384_),
    .Y(_04721_)
  );
  AND2X1 _12575_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05430_),
    .Y(_04722_)
  );
  NOR2X1 _12576_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05481_),
    .Y(_04723_)
  );
  XNOR2X1 _12577_ (
    .A(_04722_),
    .B(_04723_),
    .Y(_04724_)
  );
  NOR2X1 _12578_ (
    .A(_04721_),
    .B(_04724_),
    .Y(_04725_)
  );
  XNOR2X1 _12579_ (
    .A(_04721_),
    .B(_04724_),
    .Y(_04726_)
  );
  NOR2X1 _12580_ (
    .A(_04720_),
    .B(_04726_),
    .Y(_04727_)
  );
  XOR2X1 _12581_ (
    .A(_04720_),
    .B(_04726_),
    .Y(_04728_)
  );
  AND2X1 _12582_ (
    .A(_04719_),
    .B(_04728_),
    .Y(_04729_)
  );
  NOR2X1 _12583_ (
    .A(_04719_),
    .B(_04728_),
    .Y(_04730_)
  );
  NOR2X1 _12584_ (
    .A(_04729_),
    .B(_04730_),
    .Y(_04731_)
  );
  INVX1 _12585_ (
    .A(_04731_),
    .Y(_04732_)
  );
  NOR2X1 _12586_ (
    .A(_04712_),
    .B(_04732_),
    .Y(_04733_)
  );
  XNOR2X1 _12587_ (
    .A(_04712_),
    .B(_04731_),
    .Y(_04734_)
  );
  XOR2X1 _12588_ (
    .A(_04711_),
    .B(_04734_),
    .Y(_04735_)
  );
  XNOR2X1 _12589_ (
    .A(_04706_),
    .B(_04735_),
    .Y(_04736_)
  );
  AND2X1 _12590_ (
    .A(_04705_),
    .B(_04736_),
    .Y(_04737_)
  );
  XNOR2X1 _12591_ (
    .A(_04705_),
    .B(_04736_),
    .Y(_04738_)
  );
  AOI21X1 _12592_ (
    .A(_04684_),
    .B(_04686_),
    .C(_04738_),
    .Y(_04739_)
  );
  XNOR2X1 _12593_ (
    .A(_04703_),
    .B(_04738_),
    .Y(_04740_)
  );
  NAND2X1 _12594_ (
    .A(_04688_),
    .B(_04740_),
    .Y(_04741_)
  );
  XNOR2X1 _12595_ (
    .A(_04688_),
    .B(_04740_),
    .Y(_04742_)
  );
  XOR2X1 _12596_ (
    .A(_04702_),
    .B(_04742_),
    .Y(_04743_)
  );
  NAND2X1 _12597_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05676_),
    .Y(_04744_)
  );
  OAI21X1 _12598_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04743_),
    .C(_04744_),
    .Y(_04745_)
  );
  NAND2X1 _12599_ (
    .A(_05141_),
    .B(_04745_),
    .Y(_04746_)
  );
  NOR2X1 _12600_ (
    .A(_05141_),
    .B(_04745_),
    .Y(_04747_)
  );
  XNOR2X1 _12601_ (
    .A(multiplier_0.reshi_3_ ),
    .B(_04745_),
    .Y(_04748_)
  );
  XNOR2X1 _12602_ (
    .A(_04701_),
    .B(_04748_),
    .Y(_04749_)
  );
  AOI21X1 _12603_ (
    .A(_05225_),
    .B(_04749_),
    .C(_04590_),
    .Y(_04750_)
  );
  OAI21X1 _12604_ (
    .A(multiplier_0.reshi_3_ ),
    .B(_05225_),
    .C(_04750_),
    .Y(_04751_)
  );
  OAI21X1 _12605_ (
    .A(_05115_),
    .B(_04589_),
    .C(_04751_),
    .Y(_04440_)
  );
  OAI21X1 _12606_ (
    .A(_04702_),
    .B(_04742_),
    .C(_04741_),
    .Y(_04752_)
  );
  AOI21X1 _12607_ (
    .A(_04707_),
    .B(_04735_),
    .C(_04737_),
    .Y(_04753_)
  );
  AOI21X1 _12608_ (
    .A(_04654_),
    .B(_04710_),
    .C(_04709_),
    .Y(_04754_)
  );
  AOI21X1 _12609_ (
    .A(_04711_),
    .B(_04734_),
    .C(_04733_),
    .Y(_04755_)
  );
  OAI22X1 _12610_ (
    .A(_04664_),
    .B(_04716_),
    .C(_04718_),
    .D(_04714_),
    .Y(_04756_)
  );
  INVX1 _12611_ (
    .A(_04756_),
    .Y(_04757_)
  );
  NOR2X1 _12612_ (
    .A(_04658_),
    .B(_04757_),
    .Y(_04758_)
  );
  XNOR2X1 _12613_ (
    .A(_04658_),
    .B(_04756_),
    .Y(_04759_)
  );
  XOR2X1 _12614_ (
    .A(_04654_),
    .B(_04759_),
    .Y(_04760_)
  );
  NOR2X1 _12615_ (
    .A(_04727_),
    .B(_04729_),
    .Y(_04761_)
  );
  AOI21X1 _12616_ (
    .A(_04722_),
    .B(_04723_),
    .C(_04725_),
    .Y(_04762_)
  );
  NAND2X1 _12617_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05384_),
    .Y(_04763_)
  );
  AND2X1 _12618_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05430_),
    .Y(_04764_)
  );
  NOR2X1 _12619_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05481_),
    .Y(_04765_)
  );
  XNOR2X1 _12620_ (
    .A(_04764_),
    .B(_04765_),
    .Y(_04766_)
  );
  NOR2X1 _12621_ (
    .A(_04763_),
    .B(_04766_),
    .Y(_04767_)
  );
  XNOR2X1 _12622_ (
    .A(_04763_),
    .B(_04766_),
    .Y(_04768_)
  );
  NOR2X1 _12623_ (
    .A(_04762_),
    .B(_04768_),
    .Y(_04769_)
  );
  XOR2X1 _12624_ (
    .A(_04762_),
    .B(_04768_),
    .Y(_04770_)
  );
  OAI21X1 _12625_ (
    .A(_05302_),
    .B(_04536_),
    .C(_04716_),
    .Y(_04771_)
  );
  NAND3X1 _12626_ (
    .A(_05303_),
    .B(_05337_),
    .C(_04535_),
    .Y(_04772_)
  );
  NAND2X1 _12627_ (
    .A(_04771_),
    .B(_04772_),
    .Y(_04773_)
  );
  XNOR2X1 _12628_ (
    .A(_04713_),
    .B(_04773_),
    .Y(_04774_)
  );
  AND2X1 _12629_ (
    .A(_04770_),
    .B(_04774_),
    .Y(_04775_)
  );
  NOR2X1 _12630_ (
    .A(_04770_),
    .B(_04774_),
    .Y(_04776_)
  );
  NOR2X1 _12631_ (
    .A(_04775_),
    .B(_04776_),
    .Y(_04777_)
  );
  OAI21X1 _12632_ (
    .A(_04727_),
    .B(_04729_),
    .C(_04777_),
    .Y(_04778_)
  );
  INVX1 _12633_ (
    .A(_04778_),
    .Y(_04779_)
  );
  XNOR2X1 _12634_ (
    .A(_04761_),
    .B(_04777_),
    .Y(_04780_)
  );
  XOR2X1 _12635_ (
    .A(_04760_),
    .B(_04780_),
    .Y(_04781_)
  );
  INVX1 _12636_ (
    .A(_04781_),
    .Y(_04782_)
  );
  NOR2X1 _12637_ (
    .A(_04755_),
    .B(_04782_),
    .Y(_04783_)
  );
  XNOR2X1 _12638_ (
    .A(_04755_),
    .B(_04781_),
    .Y(_04784_)
  );
  INVX1 _12639_ (
    .A(_04784_),
    .Y(_04785_)
  );
  NOR2X1 _12640_ (
    .A(_04754_),
    .B(_04785_),
    .Y(_04786_)
  );
  XOR2X1 _12641_ (
    .A(_04754_),
    .B(_04784_),
    .Y(_04787_)
  );
  NOR2X1 _12642_ (
    .A(_04753_),
    .B(_04787_),
    .Y(_04788_)
  );
  XOR2X1 _12643_ (
    .A(_04753_),
    .B(_04787_),
    .Y(_04789_)
  );
  AND2X1 _12644_ (
    .A(_04739_),
    .B(_04789_),
    .Y(_04790_)
  );
  NOR2X1 _12645_ (
    .A(_04739_),
    .B(_04789_),
    .Y(_04791_)
  );
  NOR2X1 _12646_ (
    .A(_04790_),
    .B(_04791_),
    .Y(_04792_)
  );
  XNOR2X1 _12647_ (
    .A(_04752_),
    .B(_04792_),
    .Y(_04793_)
  );
  MUX2X1 _12648_ (
    .A(_05736_),
    .B(_04793_),
    .S(multiplier_0.cycle_0_ ),
    .Y(_04794_)
  );
  NAND2X1 _12649_ (
    .A(multiplier_0.reshi_4_ ),
    .B(_04794_),
    .Y(_04795_)
  );
  XNOR2X1 _12650_ (
    .A(multiplier_0.reshi_4_ ),
    .B(_04794_),
    .Y(_04796_)
  );
  AOI21X1 _12651_ (
    .A(_04701_),
    .B(_04746_),
    .C(_04747_),
    .Y(_04797_)
  );
  XNOR2X1 _12652_ (
    .A(_04796_),
    .B(_04797_),
    .Y(_04798_)
  );
  AOI21X1 _12653_ (
    .A(_05225_),
    .B(_04798_),
    .C(_04590_),
    .Y(_04799_)
  );
  OAI21X1 _12654_ (
    .A(multiplier_0.reshi_4_ ),
    .B(_05225_),
    .C(_04799_),
    .Y(_04800_)
  );
  OAI21X1 _12655_ (
    .A(_05117_),
    .B(_04589_),
    .C(_04800_),
    .Y(_04441_)
  );
  OAI21X1 _12656_ (
    .A(_04796_),
    .B(_04797_),
    .C(_04795_),
    .Y(_04801_)
  );
  AOI21X1 _12657_ (
    .A(_04752_),
    .B(_04792_),
    .C(_04790_),
    .Y(_04802_)
  );
  NOR2X1 _12658_ (
    .A(_04783_),
    .B(_04786_),
    .Y(_04803_)
  );
  AOI21X1 _12659_ (
    .A(_04654_),
    .B(_04759_),
    .C(_04758_),
    .Y(_04804_)
  );
  AOI21X1 _12660_ (
    .A(_04760_),
    .B(_04780_),
    .C(_04779_),
    .Y(_04805_)
  );
  OAI21X1 _12661_ (
    .A(_04714_),
    .B(_04773_),
    .C(_04772_),
    .Y(_04806_)
  );
  INVX1 _12662_ (
    .A(_04806_),
    .Y(_04807_)
  );
  NOR2X1 _12663_ (
    .A(_04658_),
    .B(_04807_),
    .Y(_04808_)
  );
  XNOR2X1 _12664_ (
    .A(_04658_),
    .B(_04806_),
    .Y(_04809_)
  );
  XNOR2X1 _12665_ (
    .A(_04654_),
    .B(_04809_),
    .Y(_04810_)
  );
  INVX1 _12666_ (
    .A(_04810_),
    .Y(_04811_)
  );
  NOR2X1 _12667_ (
    .A(_04769_),
    .B(_04775_),
    .Y(_04812_)
  );
  AOI21X1 _12668_ (
    .A(_04764_),
    .B(_04765_),
    .C(_04767_),
    .Y(_04813_)
  );
  NAND2X1 _12669_ (
    .A(multiplier_0.op1_15_ ),
    .B(_05384_),
    .Y(_04814_)
  );
  NOR2X1 _12670_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05481_),
    .Y(_04815_)
  );
  NAND3X1 _12671_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05430_),
    .C(_04815_),
    .Y(_04816_)
  );
  OAI22X1 _12672_ (
    .A(_05133_),
    .B(_05429_),
    .C(_05481_),
    .D(multiplier_0.op1_13_ ),
    .Y(_04817_)
  );
  NAND2X1 _12673_ (
    .A(_04816_),
    .B(_04817_),
    .Y(_04818_)
  );
  XNOR2X1 _12674_ (
    .A(_04814_),
    .B(_04818_),
    .Y(_04819_)
  );
  XOR2X1 _12675_ (
    .A(_04813_),
    .B(_04819_),
    .Y(_04820_)
  );
  AOI21X1 _12676_ (
    .A(_05302_),
    .B(_05336_),
    .C(_04536_),
    .Y(_04821_)
  );
  AOI22X1 _12677_ (
    .A(_04713_),
    .B(_04773_),
    .C(_04807_),
    .D(_04821_),
    .Y(_04822_)
  );
  INVX1 _12678_ (
    .A(_04822_),
    .Y(_04823_)
  );
  NAND2X1 _12679_ (
    .A(_04820_),
    .B(_04823_),
    .Y(_04824_)
  );
  XNOR2X1 _12680_ (
    .A(_04820_),
    .B(_04822_),
    .Y(_04825_)
  );
  OAI21X1 _12681_ (
    .A(_04769_),
    .B(_04775_),
    .C(_04825_),
    .Y(_04826_)
  );
  XNOR2X1 _12682_ (
    .A(_04812_),
    .B(_04825_),
    .Y(_04827_)
  );
  NAND2X1 _12683_ (
    .A(_04811_),
    .B(_04827_),
    .Y(_04828_)
  );
  XNOR2X1 _12684_ (
    .A(_04810_),
    .B(_04827_),
    .Y(_04829_)
  );
  INVX1 _12685_ (
    .A(_04829_),
    .Y(_04830_)
  );
  NOR2X1 _12686_ (
    .A(_04805_),
    .B(_04830_),
    .Y(_04831_)
  );
  XNOR2X1 _12687_ (
    .A(_04805_),
    .B(_04829_),
    .Y(_04832_)
  );
  INVX1 _12688_ (
    .A(_04832_),
    .Y(_04833_)
  );
  NOR2X1 _12689_ (
    .A(_04804_),
    .B(_04833_),
    .Y(_04834_)
  );
  XNOR2X1 _12690_ (
    .A(_04804_),
    .B(_04832_),
    .Y(_04835_)
  );
  OAI21X1 _12691_ (
    .A(_04783_),
    .B(_04786_),
    .C(_04835_),
    .Y(_04836_)
  );
  XNOR2X1 _12692_ (
    .A(_04803_),
    .B(_04835_),
    .Y(_04837_)
  );
  NAND2X1 _12693_ (
    .A(_04788_),
    .B(_04837_),
    .Y(_04838_)
  );
  XNOR2X1 _12694_ (
    .A(_04788_),
    .B(_04837_),
    .Y(_04839_)
  );
  XOR2X1 _12695_ (
    .A(_04802_),
    .B(_04839_),
    .Y(_04840_)
  );
  MUX2X1 _12696_ (
    .A(_05796_),
    .B(_04840_),
    .S(multiplier_0.cycle_0_ ),
    .Y(_04841_)
  );
  NAND2X1 _12697_ (
    .A(_05142_),
    .B(_04841_),
    .Y(_04842_)
  );
  NOR2X1 _12698_ (
    .A(_05142_),
    .B(_04841_),
    .Y(_04843_)
  );
  XNOR2X1 _12699_ (
    .A(multiplier_0.reshi_5_ ),
    .B(_04841_),
    .Y(_04844_)
  );
  XNOR2X1 _12700_ (
    .A(_04801_),
    .B(_04844_),
    .Y(_04845_)
  );
  AOI21X1 _12701_ (
    .A(_05225_),
    .B(_04845_),
    .C(_04590_),
    .Y(_04846_)
  );
  OAI21X1 _12702_ (
    .A(multiplier_0.reshi_5_ ),
    .B(_05225_),
    .C(_04846_),
    .Y(_04847_)
  );
  OAI21X1 _12703_ (
    .A(_05119_),
    .B(_04589_),
    .C(_04847_),
    .Y(_04442_)
  );
  OAI21X1 _12704_ (
    .A(_04802_),
    .B(_04839_),
    .C(_04838_),
    .Y(_04848_)
  );
  NOR2X1 _12705_ (
    .A(_04831_),
    .B(_04834_),
    .Y(_04849_)
  );
  AOI21X1 _12706_ (
    .A(_04654_),
    .B(_04809_),
    .C(_04808_),
    .Y(_04850_)
  );
  NAND2X1 _12707_ (
    .A(_04826_),
    .B(_04828_),
    .Y(_04851_)
  );
  INVX1 _12708_ (
    .A(_04851_),
    .Y(_04852_)
  );
  OAI21X1 _12709_ (
    .A(_04813_),
    .B(_04819_),
    .C(_04824_),
    .Y(_04853_)
  );
  OAI21X1 _12710_ (
    .A(_04814_),
    .B(_04818_),
    .C(_04816_),
    .Y(_04854_)
  );
  NOR2X1 _12711_ (
    .A(_05383_),
    .B(_04536_),
    .Y(_04855_)
  );
  NAND2X1 _12712_ (
    .A(multiplier_0.op1_15_ ),
    .B(_05430_),
    .Y(_04856_)
  );
  NAND2X1 _12713_ (
    .A(_05133_),
    .B(_05482_),
    .Y(_04857_)
  );
  XOR2X1 _12714_ (
    .A(_04856_),
    .B(_04857_),
    .Y(_04858_)
  );
  NAND2X1 _12715_ (
    .A(_04855_),
    .B(_04858_),
    .Y(_04859_)
  );
  XNOR2X1 _12716_ (
    .A(_04855_),
    .B(_04858_),
    .Y(_04860_)
  );
  INVX1 _12717_ (
    .A(_04860_),
    .Y(_04861_)
  );
  NAND2X1 _12718_ (
    .A(_04854_),
    .B(_04861_),
    .Y(_04862_)
  );
  XNOR2X1 _12719_ (
    .A(_04854_),
    .B(_04860_),
    .Y(_04863_)
  );
  INVX1 _12720_ (
    .A(_04863_),
    .Y(_04864_)
  );
  XNOR2X1 _12721_ (
    .A(_04822_),
    .B(_04863_),
    .Y(_04865_)
  );
  NAND2X1 _12722_ (
    .A(_04853_),
    .B(_04865_),
    .Y(_04866_)
  );
  XOR2X1 _12723_ (
    .A(_04853_),
    .B(_04865_),
    .Y(_04867_)
  );
  INVX1 _12724_ (
    .A(_04867_),
    .Y(_04868_)
  );
  XNOR2X1 _12725_ (
    .A(_04811_),
    .B(_04867_),
    .Y(_04869_)
  );
  INVX1 _12726_ (
    .A(_04869_),
    .Y(_04870_)
  );
  NOR2X1 _12727_ (
    .A(_04851_),
    .B(_04870_),
    .Y(_04871_)
  );
  XNOR2X1 _12728_ (
    .A(_04851_),
    .B(_04870_),
    .Y(_04872_)
  );
  XNOR2X1 _12729_ (
    .A(_04850_),
    .B(_04872_),
    .Y(_04873_)
  );
  NOR2X1 _12730_ (
    .A(_04849_),
    .B(_04873_),
    .Y(_04874_)
  );
  XNOR2X1 _12731_ (
    .A(_04849_),
    .B(_04873_),
    .Y(_04875_)
  );
  NOR2X1 _12732_ (
    .A(_04836_),
    .B(_04875_),
    .Y(_04876_)
  );
  XOR2X1 _12733_ (
    .A(_04836_),
    .B(_04875_),
    .Y(_04877_)
  );
  XNOR2X1 _12734_ (
    .A(_04848_),
    .B(_04877_),
    .Y(_04878_)
  );
  MUX2X1 _12735_ (
    .A(_05857_),
    .B(_04878_),
    .S(multiplier_0.cycle_0_ ),
    .Y(_04879_)
  );
  NAND2X1 _12736_ (
    .A(multiplier_0.reshi_6_ ),
    .B(_04879_),
    .Y(_04880_)
  );
  XNOR2X1 _12737_ (
    .A(multiplier_0.reshi_6_ ),
    .B(_04879_),
    .Y(_04881_)
  );
  OAI21X1 _12738_ (
    .A(_04801_),
    .B(_04843_),
    .C(_04842_),
    .Y(_04882_)
  );
  XNOR2X1 _12739_ (
    .A(_04881_),
    .B(_04882_),
    .Y(_04883_)
  );
  AOI21X1 _12740_ (
    .A(_05225_),
    .B(_04883_),
    .C(_04590_),
    .Y(_04884_)
  );
  OAI21X1 _12741_ (
    .A(multiplier_0.reshi_6_ ),
    .B(_05225_),
    .C(_04884_),
    .Y(_04885_)
  );
  OAI21X1 _12742_ (
    .A(_05121_),
    .B(_04589_),
    .C(_04885_),
    .Y(_04443_)
  );
  OAI21X1 _12743_ (
    .A(_04881_),
    .B(_04882_),
    .C(_04880_),
    .Y(_04886_)
  );
  AOI21X1 _12744_ (
    .A(_04848_),
    .B(_04877_),
    .C(_04876_),
    .Y(_04887_)
  );
  OAI21X1 _12745_ (
    .A(_04810_),
    .B(_04868_),
    .C(_04866_),
    .Y(_04888_)
  );
  OAI21X1 _12746_ (
    .A(_04822_),
    .B(_04864_),
    .C(_04862_),
    .Y(_04889_)
  );
  NAND3X1 _12747_ (
    .A(multiplier_0.op2_7_ ),
    .B(_05135_),
    .C(_04535_),
    .Y(_04890_)
  );
  OAI21X1 _12748_ (
    .A(_04856_),
    .B(_04857_),
    .C(_04859_),
    .Y(_04891_)
  );
  AOI21X1 _12749_ (
    .A(_05481_),
    .B(_04890_),
    .C(_04891_),
    .Y(_04892_)
  );
  XNOR2X1 _12750_ (
    .A(_04822_),
    .B(_04855_),
    .Y(_04893_)
  );
  XNOR2X1 _12751_ (
    .A(_04892_),
    .B(_04893_),
    .Y(_04894_)
  );
  XNOR2X1 _12752_ (
    .A(_04889_),
    .B(_04894_),
    .Y(_04895_)
  );
  XNOR2X1 _12753_ (
    .A(_04810_),
    .B(_04895_),
    .Y(_04896_)
  );
  XNOR2X1 _12754_ (
    .A(_04888_),
    .B(_04896_),
    .Y(_04897_)
  );
  OAI21X1 _12755_ (
    .A(_04852_),
    .B(_04869_),
    .C(_04850_),
    .Y(_04898_)
  );
  OAI21X1 _12756_ (
    .A(_04850_),
    .B(_04871_),
    .C(_04898_),
    .Y(_04899_)
  );
  XNOR2X1 _12757_ (
    .A(_04897_),
    .B(_04899_),
    .Y(_04900_)
  );
  XOR2X1 _12758_ (
    .A(_04874_),
    .B(_04900_),
    .Y(_04901_)
  );
  XNOR2X1 _12759_ (
    .A(_04887_),
    .B(_04901_),
    .Y(_04902_)
  );
  AND2X1 _12760_ (
    .A(_05135_),
    .B(_04902_),
    .Y(_04903_)
  );
  NOR2X1 _12761_ (
    .A(_05135_),
    .B(_04519_),
    .Y(_04904_)
  );
  NOR2X1 _12762_ (
    .A(_04903_),
    .B(_04904_),
    .Y(_04905_)
  );
  NOR2X1 _12763_ (
    .A(multiplier_0.reshi_7_ ),
    .B(_04905_),
    .Y(_04906_)
  );
  OAI21X1 _12764_ (
    .A(_04903_),
    .B(_04904_),
    .C(_05143_),
    .Y(_04907_)
  );
  NOR3X1 _12765_ (
    .A(_05143_),
    .B(_04903_),
    .C(_04904_),
    .Y(_04908_)
  );
  NOR2X1 _12766_ (
    .A(_04906_),
    .B(_04908_),
    .Y(_04909_)
  );
  XNOR2X1 _12767_ (
    .A(_04886_),
    .B(_04909_),
    .Y(_04910_)
  );
  OAI21X1 _12768_ (
    .A(multiplier_0.reshi_7_ ),
    .B(_05225_),
    .C(_04591_),
    .Y(_04911_)
  );
  AOI21X1 _12769_ (
    .A(_05225_),
    .B(_04910_),
    .C(_04911_),
    .Y(_04912_)
  );
  INVX1 _12770_ (
    .A(_04912_),
    .Y(_04913_)
  );
  OAI21X1 _12771_ (
    .A(_05123_),
    .B(_04589_),
    .C(_04913_),
    .Y(_04444_)
  );
  AOI21X1 _12772_ (
    .A(_04886_),
    .B(_04907_),
    .C(_04908_),
    .Y(_04914_)
  );
  NAND2X1 _12773_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04581_),
    .Y(_04915_)
  );
  OAI21X1 _12774_ (
    .A(_05137_),
    .B(_04902_),
    .C(_05135_),
    .Y(_04916_)
  );
  NAND2X1 _12775_ (
    .A(_04915_),
    .B(_04916_),
    .Y(_04917_)
  );
  NAND3X1 _12776_ (
    .A(multiplier_0.reshi_8_ ),
    .B(_04915_),
    .C(_04916_),
    .Y(_04918_)
  );
  AOI21X1 _12777_ (
    .A(_04915_),
    .B(_04916_),
    .C(multiplier_0.reshi_8_ ),
    .Y(_04919_)
  );
  XNOR2X1 _12778_ (
    .A(multiplier_0.reshi_8_ ),
    .B(_04917_),
    .Y(_04920_)
  );
  XNOR2X1 _12779_ (
    .A(_04914_),
    .B(_04920_),
    .Y(_04921_)
  );
  NOR2X1 _12780_ (
    .A(multiplier_0.reshi_8_ ),
    .B(_05225_),
    .Y(_04922_)
  );
  NOR2X1 _12781_ (
    .A(_04590_),
    .B(_04922_),
    .Y(_04923_)
  );
  OAI21X1 _12782_ (
    .A(_05224_),
    .B(_04921_),
    .C(_04923_),
    .Y(_04924_)
  );
  OAI21X1 _12783_ (
    .A(_05179_),
    .B(_04589_),
    .C(_04924_),
    .Y(_04445_)
  );
  OAI21X1 _12784_ (
    .A(_04914_),
    .B(_04919_),
    .C(_04918_),
    .Y(_04925_)
  );
  OAI21X1 _12785_ (
    .A(_05135_),
    .B(_04640_),
    .C(_04916_),
    .Y(_04926_)
  );
  NAND2X1 _12786_ (
    .A(_05144_),
    .B(_04926_),
    .Y(_04927_)
  );
  NOR2X1 _12787_ (
    .A(_05144_),
    .B(_04926_),
    .Y(_04928_)
  );
  XNOR2X1 _12788_ (
    .A(multiplier_0.reshi_9_ ),
    .B(_04926_),
    .Y(_04929_)
  );
  XNOR2X1 _12789_ (
    .A(_04925_),
    .B(_04929_),
    .Y(_04930_)
  );
  AOI21X1 _12790_ (
    .A(_05225_),
    .B(_04930_),
    .C(_04590_),
    .Y(_04931_)
  );
  OAI21X1 _12791_ (
    .A(multiplier_0.reshi_9_ ),
    .B(_05225_),
    .C(_04931_),
    .Y(_04932_)
  );
  OAI21X1 _12792_ (
    .A(_05181_),
    .B(_04589_),
    .C(_04932_),
    .Y(_04446_)
  );
  NAND2X1 _12793_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04693_),
    .Y(_04933_)
  );
  NAND2X1 _12794_ (
    .A(_04916_),
    .B(_04933_),
    .Y(_04934_)
  );
  NAND3X1 _12795_ (
    .A(multiplier_0.reshi_10_ ),
    .B(_04916_),
    .C(_04933_),
    .Y(_04935_)
  );
  XOR2X1 _12796_ (
    .A(multiplier_0.reshi_10_ ),
    .B(_04934_),
    .Y(_04936_)
  );
  AOI21X1 _12797_ (
    .A(_04925_),
    .B(_04927_),
    .C(_04928_),
    .Y(_04937_)
  );
  XNOR2X1 _12798_ (
    .A(_04936_),
    .B(_04937_),
    .Y(_04938_)
  );
  AOI21X1 _12799_ (
    .A(_05225_),
    .B(_04938_),
    .C(_04590_),
    .Y(_04939_)
  );
  OAI21X1 _12800_ (
    .A(multiplier_0.reshi_10_ ),
    .B(_05225_),
    .C(_04939_),
    .Y(_04940_)
  );
  OAI21X1 _12801_ (
    .A(_05183_),
    .B(_04589_),
    .C(_04940_),
    .Y(_04432_)
  );
  OAI21X1 _12802_ (
    .A(_04936_),
    .B(_04937_),
    .C(_04935_),
    .Y(_04941_)
  );
  OAI21X1 _12803_ (
    .A(_05135_),
    .B(_04743_),
    .C(_04916_),
    .Y(_04942_)
  );
  NAND2X1 _12804_ (
    .A(_05145_),
    .B(_04942_),
    .Y(_04943_)
  );
  NOR2X1 _12805_ (
    .A(_05145_),
    .B(_04942_),
    .Y(_04944_)
  );
  XNOR2X1 _12806_ (
    .A(multiplier_0.reshi_11_ ),
    .B(_04942_),
    .Y(_04945_)
  );
  XNOR2X1 _12807_ (
    .A(_04941_),
    .B(_04945_),
    .Y(_04946_)
  );
  AOI21X1 _12808_ (
    .A(_05225_),
    .B(_04946_),
    .C(_04590_),
    .Y(_04947_)
  );
  OAI21X1 _12809_ (
    .A(multiplier_0.reshi_11_ ),
    .B(_05225_),
    .C(_04947_),
    .Y(_04948_)
  );
  OAI21X1 _12810_ (
    .A(_05185_),
    .B(_04589_),
    .C(_04948_),
    .Y(_04433_)
  );
  NAND2X1 _12811_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04793_),
    .Y(_04949_)
  );
  NAND2X1 _12812_ (
    .A(_04916_),
    .B(_04949_),
    .Y(_04950_)
  );
  NAND3X1 _12813_ (
    .A(multiplier_0.reshi_12_ ),
    .B(_04916_),
    .C(_04949_),
    .Y(_04951_)
  );
  XOR2X1 _12814_ (
    .A(multiplier_0.reshi_12_ ),
    .B(_04950_),
    .Y(_04952_)
  );
  AOI21X1 _12815_ (
    .A(_04941_),
    .B(_04943_),
    .C(_04944_),
    .Y(_04953_)
  );
  XOR2X1 _12816_ (
    .A(_04952_),
    .B(_04953_),
    .Y(_04954_)
  );
  NOR2X1 _12817_ (
    .A(multiplier_0.reshi_12_ ),
    .B(_05225_),
    .Y(_04955_)
  );
  NOR2X1 _12818_ (
    .A(_04590_),
    .B(_04955_),
    .Y(_04956_)
  );
  OAI21X1 _12819_ (
    .A(_05224_),
    .B(_04954_),
    .C(_04956_),
    .Y(_04957_)
  );
  OAI21X1 _12820_ (
    .A(_05187_),
    .B(_04589_),
    .C(_04957_),
    .Y(_04434_)
  );
  OAI21X1 _12821_ (
    .A(_04952_),
    .B(_04953_),
    .C(_04951_),
    .Y(_04958_)
  );
  OAI21X1 _12822_ (
    .A(_05135_),
    .B(_04840_),
    .C(_04916_),
    .Y(_04959_)
  );
  NAND2X1 _12823_ (
    .A(_05146_),
    .B(_04959_),
    .Y(_04960_)
  );
  NOR2X1 _12824_ (
    .A(_05146_),
    .B(_04959_),
    .Y(_04961_)
  );
  XNOR2X1 _12825_ (
    .A(multiplier_0.reshi_13_ ),
    .B(_04959_),
    .Y(_04962_)
  );
  XNOR2X1 _12826_ (
    .A(_04958_),
    .B(_04962_),
    .Y(_04963_)
  );
  AOI21X1 _12827_ (
    .A(_05225_),
    .B(_04963_),
    .C(_04590_),
    .Y(_04964_)
  );
  OAI21X1 _12828_ (
    .A(multiplier_0.reshi_13_ ),
    .B(_05225_),
    .C(_04964_),
    .Y(_04965_)
  );
  OAI21X1 _12829_ (
    .A(_05189_),
    .B(_04589_),
    .C(_04965_),
    .Y(_04435_)
  );
  NAND2X1 _12830_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04878_),
    .Y(_04966_)
  );
  NAND2X1 _12831_ (
    .A(_04916_),
    .B(_04966_),
    .Y(_04967_)
  );
  NAND3X1 _12832_ (
    .A(multiplier_0.reshi_14_ ),
    .B(_04916_),
    .C(_04966_),
    .Y(_04968_)
  );
  XOR2X1 _12833_ (
    .A(multiplier_0.reshi_14_ ),
    .B(_04967_),
    .Y(_04969_)
  );
  OAI21X1 _12834_ (
    .A(_04958_),
    .B(_04961_),
    .C(_04960_),
    .Y(_04970_)
  );
  XNOR2X1 _12835_ (
    .A(_04969_),
    .B(_04970_),
    .Y(_04971_)
  );
  AOI21X1 _12836_ (
    .A(_05225_),
    .B(_04971_),
    .C(_04590_),
    .Y(_04972_)
  );
  OAI21X1 _12837_ (
    .A(multiplier_0.reshi_14_ ),
    .B(_05225_),
    .C(_04972_),
    .Y(_04973_)
  );
  OAI21X1 _12838_ (
    .A(_05191_),
    .B(_04589_),
    .C(_04973_),
    .Y(_04436_)
  );
  OAI21X1 _12839_ (
    .A(_04969_),
    .B(_04970_),
    .C(_04968_),
    .Y(_04974_)
  );
  AOI21X1 _12840_ (
    .A(_05135_),
    .B(_05137_),
    .C(_04902_),
    .Y(_04975_)
  );
  XOR2X1 _12841_ (
    .A(multiplier_0.reshi_15_ ),
    .B(_04975_),
    .Y(_04976_)
  );
  NAND2X1 _12842_ (
    .A(_04974_),
    .B(_04976_),
    .Y(_04977_)
  );
  XNOR2X1 _12843_ (
    .A(_04974_),
    .B(_04976_),
    .Y(_04978_)
  );
  AOI21X1 _12844_ (
    .A(_05225_),
    .B(_04978_),
    .C(_04590_),
    .Y(_04979_)
  );
  OAI21X1 _12845_ (
    .A(multiplier_0.reshi_15_ ),
    .B(_05225_),
    .C(_04979_),
    .Y(_04980_)
  );
  OAI21X1 _12846_ (
    .A(_05193_),
    .B(_04589_),
    .C(_04980_),
    .Y(_04437_)
  );
  NOR2X1 _12847_ (
    .A(_05137_),
    .B(_04978_),
    .Y(_04981_)
  );
  AOI21X1 _12848_ (
    .A(multiplier_0.reshi_15_ ),
    .B(_04975_),
    .C(multiplier_0.sumext_0_ ),
    .Y(_04982_)
  );
  AOI21X1 _12849_ (
    .A(_04977_),
    .B(_04982_),
    .C(multiplier_0.sign_sel ),
    .Y(_04983_)
  );
  NOR2X1 _12850_ (
    .A(_04981_),
    .B(_04983_),
    .Y(_04984_)
  );
  OAI21X1 _12851_ (
    .A(multiplier_0.sumext_0_ ),
    .B(_05225_),
    .C(_05169_),
    .Y(_04985_)
  );
  AOI21X1 _12852_ (
    .A(_05225_),
    .B(_04984_),
    .C(_04985_),
    .Y(_04464_)
  );
  NOR2X1 _12853_ (
    .A(_05224_),
    .B(_04981_),
    .Y(_04986_)
  );
  OAI21X1 _12854_ (
    .A(multiplier_0.sumext_10_ ),
    .B(_05225_),
    .C(_05161_),
    .Y(_04987_)
  );
  NOR2X1 _12855_ (
    .A(_04986_),
    .B(_04987_),
    .Y(_04465_)
  );
  MUX2X1 _12856_ (
    .A(multiplier_0.acc_sel ),
    .B(_00101_),
    .S(_05194_),
    .Y(_04988_)
  );
  INVX1 _12857_ (
    .A(_04988_),
    .Y(_04398_)
  );
  MUX2X1 _12858_ (
    .A(multiplier_0.sign_sel ),
    .B(_00097_),
    .S(_05194_),
    .Y(_04989_)
  );
  INVX1 _12859_ (
    .A(_04989_),
    .Y(_04463_)
  );
  NOR3X1 _12860_ (
    .A(_05136_),
    .B(_04981_),
    .C(_04983_),
    .Y(_04990_)
  );
  NAND2X1 _12861_ (
    .A(_05156_),
    .B(_05157_),
    .Y(_04991_)
  );
  NAND3X1 _12862_ (
    .A(_00101_),
    .B(_05156_),
    .C(_05157_),
    .Y(_04992_)
  );
  NOR2X1 _12863_ (
    .A(_05217_),
    .B(_04992_),
    .Y(_04993_)
  );
  OAI21X1 _12864_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.sumext_0_ ),
    .C(_04993_),
    .Y(_04994_)
  );
  NOR2X1 _12865_ (
    .A(_05136_),
    .B(_04586_),
    .Y(_04995_)
  );
  NOR2X1 _12866_ (
    .A(_05159_),
    .B(_04992_),
    .Y(_04996_)
  );
  OAI21X1 _12867_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_0_ ),
    .C(_04996_),
    .Y(_04997_)
  );
  NOR2X1 _12868_ (
    .A(_04995_),
    .B(_04997_),
    .Y(_04998_)
  );
  NOR2X1 _12869_ (
    .A(_05160_),
    .B(_04991_),
    .Y(_04999_)
  );
  NAND2X1 _12870_ (
    .A(multiplier_0.op2_0_ ),
    .B(_04999_),
    .Y(_05000_)
  );
  NOR2X1 _12871_ (
    .A(_05218_),
    .B(_04991_),
    .Y(_05001_)
  );
  OR2X1 _12872_ (
    .A(_05218_),
    .B(_04991_),
    .Y(_05002_)
  );
  NOR2X1 _12873_ (
    .A(_00102_),
    .B(_04991_),
    .Y(_05003_)
  );
  AOI22X1 _12874_ (
    .A(_05216_),
    .B(_05001_),
    .C(_05003_),
    .D(multiplier_0.op1_0_ ),
    .Y(_05004_)
  );
  NAND2X1 _12875_ (
    .A(_05000_),
    .B(_05004_),
    .Y(_05005_)
  );
  NOR2X1 _12876_ (
    .A(_04998_),
    .B(_05005_),
    .Y(_05006_)
  );
  OAI21X1 _12877_ (
    .A(_04990_),
    .B(_04994_),
    .C(_05006_),
    .Y(multiplier_0.per_dout_0_ )
  );
  OAI21X1 _12878_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.sumext_10_ ),
    .C(_04993_),
    .Y(_05007_)
  );
  INVX1 _12879_ (
    .A(_05007_),
    .Y(_05008_)
  );
  OAI21X1 _12880_ (
    .A(_05136_),
    .B(_04981_),
    .C(_05008_),
    .Y(_05009_)
  );
  OAI21X1 _12881_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_1_ ),
    .C(_04996_),
    .Y(_05010_)
  );
  AOI21X1 _12882_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04646_),
    .C(_05010_),
    .Y(_05011_)
  );
  AOI22X1 _12883_ (
    .A(multiplier_0.op2_1_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_1_ ),
    .Y(_05012_)
  );
  OAI21X1 _12884_ (
    .A(_05240_),
    .B(_05002_),
    .C(_05012_),
    .Y(_05013_)
  );
  NOR2X1 _12885_ (
    .A(_05011_),
    .B(_05013_),
    .Y(_05014_)
  );
  NAND2X1 _12886_ (
    .A(_05009_),
    .B(_05014_),
    .Y(multiplier_0.per_dout_1_ )
  );
  OAI21X1 _12887_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_2_ ),
    .C(_04996_),
    .Y(_05015_)
  );
  AOI21X1 _12888_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04698_),
    .C(_05015_),
    .Y(_05016_)
  );
  AOI22X1 _12889_ (
    .A(multiplier_0.op2_2_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_2_ ),
    .Y(_05017_)
  );
  OAI21X1 _12890_ (
    .A(_05260_),
    .B(_05002_),
    .C(_05017_),
    .Y(_05018_)
  );
  NOR2X1 _12891_ (
    .A(_05016_),
    .B(_05018_),
    .Y(_05019_)
  );
  NAND2X1 _12892_ (
    .A(_05009_),
    .B(_05019_),
    .Y(multiplier_0.per_dout_2_ )
  );
  OAI21X1 _12893_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_3_ ),
    .C(_04996_),
    .Y(_05020_)
  );
  AOI21X1 _12894_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04749_),
    .C(_05020_),
    .Y(_05021_)
  );
  AOI22X1 _12895_ (
    .A(multiplier_0.op2_3_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_3_ ),
    .Y(_05022_)
  );
  OAI21X1 _12896_ (
    .A(_05288_),
    .B(_05002_),
    .C(_05022_),
    .Y(_05023_)
  );
  NOR2X1 _12897_ (
    .A(_05021_),
    .B(_05023_),
    .Y(_05024_)
  );
  NAND2X1 _12898_ (
    .A(_05009_),
    .B(_05024_),
    .Y(multiplier_0.per_dout_3_ )
  );
  OAI21X1 _12899_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_4_ ),
    .C(_04996_),
    .Y(_05025_)
  );
  AOI21X1 _12900_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04798_),
    .C(_05025_),
    .Y(_05026_)
  );
  AOI22X1 _12901_ (
    .A(multiplier_0.op2_4_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_4_ ),
    .Y(_05027_)
  );
  OAI21X1 _12902_ (
    .A(_05320_),
    .B(_05002_),
    .C(_05027_),
    .Y(_05028_)
  );
  NOR2X1 _12903_ (
    .A(_05026_),
    .B(_05028_),
    .Y(_05029_)
  );
  NAND2X1 _12904_ (
    .A(_05009_),
    .B(_05029_),
    .Y(multiplier_0.per_dout_4_ )
  );
  OAI21X1 _12905_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_5_ ),
    .C(_04996_),
    .Y(_05030_)
  );
  AOI21X1 _12906_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04845_),
    .C(_05030_),
    .Y(_05031_)
  );
  AOI22X1 _12907_ (
    .A(multiplier_0.op2_5_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_5_ ),
    .Y(_05032_)
  );
  OAI21X1 _12908_ (
    .A(_05359_),
    .B(_05002_),
    .C(_05032_),
    .Y(_05033_)
  );
  NOR2X1 _12909_ (
    .A(_05031_),
    .B(_05033_),
    .Y(_05034_)
  );
  NAND2X1 _12910_ (
    .A(_05009_),
    .B(_05034_),
    .Y(multiplier_0.per_dout_5_ )
  );
  OAI21X1 _12911_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_6_ ),
    .C(_04996_),
    .Y(_05035_)
  );
  AOI21X1 _12912_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04883_),
    .C(_05035_),
    .Y(_05036_)
  );
  AOI22X1 _12913_ (
    .A(multiplier_0.op2_6_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_6_ ),
    .Y(_05037_)
  );
  OAI21X1 _12914_ (
    .A(_05403_),
    .B(_05002_),
    .C(_05037_),
    .Y(_05038_)
  );
  NOR2X1 _12915_ (
    .A(_05036_),
    .B(_05038_),
    .Y(_05039_)
  );
  NAND2X1 _12916_ (
    .A(_05009_),
    .B(_05039_),
    .Y(multiplier_0.per_dout_6_ )
  );
  OAI21X1 _12917_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_7_ ),
    .C(_04996_),
    .Y(_05040_)
  );
  AOI21X1 _12918_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04910_),
    .C(_05040_),
    .Y(_05041_)
  );
  AOI22X1 _12919_ (
    .A(multiplier_0.op2_7_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_7_ ),
    .Y(_05042_)
  );
  OAI21X1 _12920_ (
    .A(_05454_),
    .B(_05002_),
    .C(_05042_),
    .Y(_05043_)
  );
  NOR2X1 _12921_ (
    .A(_05041_),
    .B(_05043_),
    .Y(_05044_)
  );
  NAND2X1 _12922_ (
    .A(_05009_),
    .B(_05044_),
    .Y(multiplier_0.per_dout_7_ )
  );
  NOR2X1 _12923_ (
    .A(_05136_),
    .B(_04921_),
    .Y(_05045_)
  );
  OAI21X1 _12924_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_8_ ),
    .C(_04996_),
    .Y(_05046_)
  );
  NOR2X1 _12925_ (
    .A(_05045_),
    .B(_05046_),
    .Y(_05047_)
  );
  NOR2X1 _12926_ (
    .A(_05136_),
    .B(_05507_),
    .Y(_05048_)
  );
  OAI21X1 _12927_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_8_ ),
    .C(_05001_),
    .Y(_05049_)
  );
  AOI22X1 _12928_ (
    .A(multiplier_0.op2_8_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_8_ ),
    .Y(_05050_)
  );
  OAI21X1 _12929_ (
    .A(_05048_),
    .B(_05049_),
    .C(_05050_),
    .Y(_05051_)
  );
  NOR2X1 _12930_ (
    .A(_05047_),
    .B(_05051_),
    .Y(_05052_)
  );
  NAND2X1 _12931_ (
    .A(_05009_),
    .B(_05052_),
    .Y(multiplier_0.per_dout_8_ )
  );
  OAI21X1 _12932_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_9_ ),
    .C(_04996_),
    .Y(_05053_)
  );
  AOI21X1 _12933_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04930_),
    .C(_05053_),
    .Y(_05054_)
  );
  NOR2X1 _12934_ (
    .A(_05136_),
    .B(_05566_),
    .Y(_05055_)
  );
  OAI21X1 _12935_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_9_ ),
    .C(_05001_),
    .Y(_05056_)
  );
  AOI22X1 _12936_ (
    .A(multiplier_0.op2_9_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_9_ ),
    .Y(_05057_)
  );
  OAI21X1 _12937_ (
    .A(_05055_),
    .B(_05056_),
    .C(_05057_),
    .Y(_05058_)
  );
  NOR2X1 _12938_ (
    .A(_05054_),
    .B(_05058_),
    .Y(_05059_)
  );
  NAND2X1 _12939_ (
    .A(_05009_),
    .B(_05059_),
    .Y(multiplier_0.per_dout_9_ )
  );
  OAI21X1 _12940_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_10_ ),
    .C(_04996_),
    .Y(_05060_)
  );
  AOI21X1 _12941_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04938_),
    .C(_05060_),
    .Y(_05061_)
  );
  AND2X1 _12942_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_05622_),
    .Y(_05062_)
  );
  OAI21X1 _12943_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_10_ ),
    .C(_05001_),
    .Y(_05063_)
  );
  AOI22X1 _12944_ (
    .A(multiplier_0.op2_10_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_10_ ),
    .Y(_05064_)
  );
  OAI21X1 _12945_ (
    .A(_05062_),
    .B(_05063_),
    .C(_05064_),
    .Y(_05065_)
  );
  NOR2X1 _12946_ (
    .A(_05061_),
    .B(_05065_),
    .Y(_05066_)
  );
  NAND2X1 _12947_ (
    .A(_05009_),
    .B(_05066_),
    .Y(multiplier_0.per_dout_10_ )
  );
  OAI21X1 _12948_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_11_ ),
    .C(_04996_),
    .Y(_05067_)
  );
  AOI21X1 _12949_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04946_),
    .C(_05067_),
    .Y(_05068_)
  );
  AND2X1 _12950_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_05680_),
    .Y(_05069_)
  );
  OAI21X1 _12951_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_11_ ),
    .C(_05001_),
    .Y(_05070_)
  );
  AOI22X1 _12952_ (
    .A(multiplier_0.op2_11_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_11_ ),
    .Y(_05071_)
  );
  OAI21X1 _12953_ (
    .A(_05069_),
    .B(_05070_),
    .C(_05071_),
    .Y(_05072_)
  );
  NOR2X1 _12954_ (
    .A(_05068_),
    .B(_05072_),
    .Y(_05073_)
  );
  NAND2X1 _12955_ (
    .A(_05009_),
    .B(_05073_),
    .Y(multiplier_0.per_dout_11_ )
  );
  NOR2X1 _12956_ (
    .A(_05136_),
    .B(_04954_),
    .Y(_05074_)
  );
  OAI21X1 _12957_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_12_ ),
    .C(_04996_),
    .Y(_05075_)
  );
  NOR2X1 _12958_ (
    .A(_05074_),
    .B(_05075_),
    .Y(_05076_)
  );
  NOR2X1 _12959_ (
    .A(_05136_),
    .B(_05741_),
    .Y(_05077_)
  );
  OAI21X1 _12960_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_12_ ),
    .C(_05001_),
    .Y(_05078_)
  );
  AOI22X1 _12961_ (
    .A(multiplier_0.op2_12_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_12_ ),
    .Y(_05079_)
  );
  OAI21X1 _12962_ (
    .A(_05077_),
    .B(_05078_),
    .C(_05079_),
    .Y(_05080_)
  );
  NOR2X1 _12963_ (
    .A(_05076_),
    .B(_05080_),
    .Y(_05081_)
  );
  NAND2X1 _12964_ (
    .A(_05009_),
    .B(_05081_),
    .Y(multiplier_0.per_dout_12_ )
  );
  OAI21X1 _12965_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_13_ ),
    .C(_04996_),
    .Y(_05082_)
  );
  AOI21X1 _12966_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04963_),
    .C(_05082_),
    .Y(_05083_)
  );
  AND2X1 _12967_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_05801_),
    .Y(_05084_)
  );
  OAI21X1 _12968_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_13_ ),
    .C(_05001_),
    .Y(_05085_)
  );
  AOI22X1 _12969_ (
    .A(multiplier_0.op2_13_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_13_ ),
    .Y(_05086_)
  );
  OAI21X1 _12970_ (
    .A(_05084_),
    .B(_05085_),
    .C(_05086_),
    .Y(_05087_)
  );
  NOR2X1 _12971_ (
    .A(_05083_),
    .B(_05087_),
    .Y(_05088_)
  );
  NAND2X1 _12972_ (
    .A(_05009_),
    .B(_05088_),
    .Y(multiplier_0.per_dout_13_ )
  );
  OAI21X1 _12973_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_14_ ),
    .C(_04996_),
    .Y(_05089_)
  );
  AOI21X1 _12974_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04971_),
    .C(_05089_),
    .Y(_05090_)
  );
  NOR2X1 _12975_ (
    .A(_05136_),
    .B(_05863_),
    .Y(_05091_)
  );
  OAI21X1 _12976_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_14_ ),
    .C(_05001_),
    .Y(_05092_)
  );
  AOI22X1 _12977_ (
    .A(multiplier_0.op2_14_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_14_ ),
    .Y(_05093_)
  );
  OAI21X1 _12978_ (
    .A(_05091_),
    .B(_05092_),
    .C(_05093_),
    .Y(_05094_)
  );
  NOR2X1 _12979_ (
    .A(_05090_),
    .B(_05094_),
    .Y(_05095_)
  );
  NAND2X1 _12980_ (
    .A(_05009_),
    .B(_05095_),
    .Y(multiplier_0.per_dout_14_ )
  );
  OAI21X1 _12981_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_15_ ),
    .C(_04996_),
    .Y(_05096_)
  );
  AOI21X1 _12982_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04978_),
    .C(_05096_),
    .Y(_05097_)
  );
  AND2X1 _12983_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04524_),
    .Y(_05098_)
  );
  OAI21X1 _12984_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_15_ ),
    .C(_05001_),
    .Y(_05099_)
  );
  AOI22X1 _12985_ (
    .A(multiplier_0.op2_15_ ),
    .B(_04999_),
    .C(_05003_),
    .D(multiplier_0.op1_15_ ),
    .Y(_05100_)
  );
  OAI21X1 _12986_ (
    .A(_05098_),
    .B(_05099_),
    .C(_05100_),
    .Y(_05101_)
  );
  NOR2X1 _12987_ (
    .A(_05097_),
    .B(_05101_),
    .Y(_05102_)
  );
  NAND2X1 _12988_ (
    .A(_05009_),
    .B(_05102_),
    .Y(multiplier_0.per_dout_15_ )
  );
  DFFSR _12989_ (
    .CLK(dco_clk),
    .D(multiplier_0.op2_wr ),
    .Q(multiplier_0.cycle_0_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _12990_ (
    .CLK(dco_clk),
    .D(multiplier_0.cycle_0_ ),
    .Q(multiplier_0.cycle_1_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _12991_ (
    .CLK(dco_clk),
    .D(_04398_),
    .Q(multiplier_0.acc_sel ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _12992_ (
    .CLK(dco_clk),
    .D(_04463_),
    .Q(multiplier_0.sign_sel ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _12993_ (
    .CLK(dco_clk),
    .D(_04464_),
    .Q(multiplier_0.sumext_0_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _12994_ (
    .CLK(dco_clk),
    .D(_04465_),
    .Q(multiplier_0.sumext_10_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _12995_ (
    .CLK(dco_clk),
    .D(_04431_),
    .Q(multiplier_0.reshi_0_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _12996_ (
    .CLK(dco_clk),
    .D(_04438_),
    .Q(multiplier_0.reshi_1_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _12997_ (
    .CLK(dco_clk),
    .D(_04439_),
    .Q(multiplier_0.reshi_2_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _12998_ (
    .CLK(dco_clk),
    .D(_04440_),
    .Q(multiplier_0.reshi_3_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _12999_ (
    .CLK(dco_clk),
    .D(_04441_),
    .Q(multiplier_0.reshi_4_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13000_ (
    .CLK(dco_clk),
    .D(_04442_),
    .Q(multiplier_0.reshi_5_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13001_ (
    .CLK(dco_clk),
    .D(_04443_),
    .Q(multiplier_0.reshi_6_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13002_ (
    .CLK(dco_clk),
    .D(_04444_),
    .Q(multiplier_0.reshi_7_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13003_ (
    .CLK(dco_clk),
    .D(_04445_),
    .Q(multiplier_0.reshi_8_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13004_ (
    .CLK(dco_clk),
    .D(_04446_),
    .Q(multiplier_0.reshi_9_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13005_ (
    .CLK(dco_clk),
    .D(_04432_),
    .Q(multiplier_0.reshi_10_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13006_ (
    .CLK(dco_clk),
    .D(_04433_),
    .Q(multiplier_0.reshi_11_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13007_ (
    .CLK(dco_clk),
    .D(_04434_),
    .Q(multiplier_0.reshi_12_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13008_ (
    .CLK(dco_clk),
    .D(_04435_),
    .Q(multiplier_0.reshi_13_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13009_ (
    .CLK(dco_clk),
    .D(_04436_),
    .Q(multiplier_0.reshi_14_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13010_ (
    .CLK(dco_clk),
    .D(_04437_),
    .Q(multiplier_0.reshi_15_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13011_ (
    .CLK(dco_clk),
    .D(_04447_),
    .Q(multiplier_0.reslo_0_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13012_ (
    .CLK(dco_clk),
    .D(_04454_),
    .Q(multiplier_0.reslo_1_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13013_ (
    .CLK(dco_clk),
    .D(_04455_),
    .Q(multiplier_0.reslo_2_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13014_ (
    .CLK(dco_clk),
    .D(_04456_),
    .Q(multiplier_0.reslo_3_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13015_ (
    .CLK(dco_clk),
    .D(_04457_),
    .Q(multiplier_0.reslo_4_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13016_ (
    .CLK(dco_clk),
    .D(_04458_),
    .Q(multiplier_0.reslo_5_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13017_ (
    .CLK(dco_clk),
    .D(_04459_),
    .Q(multiplier_0.reslo_6_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13018_ (
    .CLK(dco_clk),
    .D(_04460_),
    .Q(multiplier_0.reslo_7_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13019_ (
    .CLK(dco_clk),
    .D(_04461_),
    .Q(multiplier_0.reslo_8_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13020_ (
    .CLK(dco_clk),
    .D(_04462_),
    .Q(multiplier_0.reslo_9_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13021_ (
    .CLK(dco_clk),
    .D(_04448_),
    .Q(multiplier_0.reslo_10_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13022_ (
    .CLK(dco_clk),
    .D(_04449_),
    .Q(multiplier_0.reslo_11_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13023_ (
    .CLK(dco_clk),
    .D(_04450_),
    .Q(multiplier_0.reslo_12_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13024_ (
    .CLK(dco_clk),
    .D(_04451_),
    .Q(multiplier_0.reslo_13_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13025_ (
    .CLK(dco_clk),
    .D(_04452_),
    .Q(multiplier_0.reslo_14_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13026_ (
    .CLK(dco_clk),
    .D(_04453_),
    .Q(multiplier_0.reslo_15_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13027_ (
    .CLK(dco_clk),
    .D(_04415_),
    .Q(multiplier_0.op2_0_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13028_ (
    .CLK(dco_clk),
    .D(_04422_),
    .Q(multiplier_0.op2_1_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13029_ (
    .CLK(dco_clk),
    .D(_04423_),
    .Q(multiplier_0.op2_2_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13030_ (
    .CLK(dco_clk),
    .D(_04424_),
    .Q(multiplier_0.op2_3_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13031_ (
    .CLK(dco_clk),
    .D(_04425_),
    .Q(multiplier_0.op2_4_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13032_ (
    .CLK(dco_clk),
    .D(_04426_),
    .Q(multiplier_0.op2_5_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13033_ (
    .CLK(dco_clk),
    .D(_04427_),
    .Q(multiplier_0.op2_6_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13034_ (
    .CLK(dco_clk),
    .D(_04428_),
    .Q(multiplier_0.op2_7_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13035_ (
    .CLK(dco_clk),
    .D(_04429_),
    .Q(multiplier_0.op2_8_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13036_ (
    .CLK(dco_clk),
    .D(_04430_),
    .Q(multiplier_0.op2_9_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13037_ (
    .CLK(dco_clk),
    .D(_04416_),
    .Q(multiplier_0.op2_10_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13038_ (
    .CLK(dco_clk),
    .D(_04417_),
    .Q(multiplier_0.op2_11_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13039_ (
    .CLK(dco_clk),
    .D(_04418_),
    .Q(multiplier_0.op2_12_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13040_ (
    .CLK(dco_clk),
    .D(_04419_),
    .Q(multiplier_0.op2_13_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13041_ (
    .CLK(dco_clk),
    .D(_04420_),
    .Q(multiplier_0.op2_14_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13042_ (
    .CLK(dco_clk),
    .D(_04421_),
    .Q(multiplier_0.op2_15_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13043_ (
    .CLK(dco_clk),
    .D(_04399_),
    .Q(multiplier_0.op1_0_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13044_ (
    .CLK(dco_clk),
    .D(_04406_),
    .Q(multiplier_0.op1_1_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13045_ (
    .CLK(dco_clk),
    .D(_04407_),
    .Q(multiplier_0.op1_2_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13046_ (
    .CLK(dco_clk),
    .D(_04408_),
    .Q(multiplier_0.op1_3_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13047_ (
    .CLK(dco_clk),
    .D(_04409_),
    .Q(multiplier_0.op1_4_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13048_ (
    .CLK(dco_clk),
    .D(_04410_),
    .Q(multiplier_0.op1_5_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13049_ (
    .CLK(dco_clk),
    .D(_04411_),
    .Q(multiplier_0.op1_6_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13050_ (
    .CLK(dco_clk),
    .D(_04412_),
    .Q(multiplier_0.op1_7_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13051_ (
    .CLK(dco_clk),
    .D(_04413_),
    .Q(multiplier_0.op1_8_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13052_ (
    .CLK(dco_clk),
    .D(_04414_),
    .Q(multiplier_0.op1_9_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13053_ (
    .CLK(dco_clk),
    .D(_04400_),
    .Q(multiplier_0.op1_10_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13054_ (
    .CLK(dco_clk),
    .D(_04401_),
    .Q(multiplier_0.op1_11_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13055_ (
    .CLK(dco_clk),
    .D(_04402_),
    .Q(multiplier_0.op1_12_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13056_ (
    .CLK(dco_clk),
    .D(_04403_),
    .Q(multiplier_0.op1_13_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13057_ (
    .CLK(dco_clk),
    .D(_04404_),
    .Q(multiplier_0.op1_14_ ),
    .R(_04466_),
    .S(1'h1)
  );
  DFFSR _13058_ (
    .CLK(dco_clk),
    .D(_04405_),
    .Q(multiplier_0.op1_15_ ),
    .R(_04466_),
    .S(1'h1)
  );
  INVX1 _13059_ (
    .A(_00101_),
    .Y(_05874_)
  );
  INVX1 _13060_ (
    .A(_00102_),
    .Y(_05875_)
  );
  INVX1 _13061_ (
    .A(_00100_),
    .Y(_05876_)
  );
  INVX1 _13062_ (
    .A(_00126_),
    .Y(_05877_)
  );
  INVX1 _13063_ (
    .A(_00110_),
    .Y(_05878_)
  );
  INVX1 _13064_ (
    .A(sfr_0.ie1_0_ ),
    .Y(_05879_)
  );
  INVX1 _13065_ (
    .A(1'h0),
    .Y(_05880_)
  );
  INVX1 _13066_ (
    .A(1'h0),
    .Y(_05881_)
  );
  INVX1 _13067_ (
    .A(1'h0),
    .Y(_05882_)
  );
  INVX1 _13068_ (
    .A(1'h0),
    .Y(_05883_)
  );
  INVX1 _13069_ (
    .A(sfr_0.ifg1_0_ ),
    .Y(_05884_)
  );
  INVX1 _13070_ (
    .A(_00162_),
    .Y(_05865_)
  );
  NOR2X1 _13071_ (
    .A(_00097_),
    .B(_00101_),
    .Y(_05885_)
  );
  AND2X1 _13072_ (
    .A(_05875_),
    .B(_05885_),
    .Y(_05886_)
  );
  NOR2X1 _13073_ (
    .A(_00099_),
    .B(1'h0),
    .Y(_05887_)
  );
  OR2X1 _13074_ (
    .A(_00099_),
    .B(1'h0),
    .Y(_05888_)
  );
  NOR3X1 _13075_ (
    .A(_00100_),
    .B(_05877_),
    .C(_05888_),
    .Y(_05889_)
  );
  NAND3X1 _13076_ (
    .A(_05876_),
    .B(_00126_),
    .C(_05887_),
    .Y(_05890_)
  );
  NOR2X1 _13077_ (
    .A(_00108_),
    .B(_00107_),
    .Y(_05891_)
  );
  NOR2X1 _13078_ (
    .A(_00098_),
    .B(_00109_),
    .Y(_05892_)
  );
  AND2X1 _13079_ (
    .A(_05891_),
    .B(_05892_),
    .Y(_05893_)
  );
  NAND2X1 _13080_ (
    .A(_05891_),
    .B(_05892_),
    .Y(_05894_)
  );
  NOR2X1 _13081_ (
    .A(_00104_),
    .B(_00103_),
    .Y(_05895_)
  );
  NOR2X1 _13082_ (
    .A(_00106_),
    .B(_00105_),
    .Y(_05896_)
  );
  AND2X1 _13083_ (
    .A(_05895_),
    .B(_05896_),
    .Y(_05897_)
  );
  NAND2X1 _13084_ (
    .A(_05895_),
    .B(_05896_),
    .Y(_05898_)
  );
  NOR3X1 _13085_ (
    .A(_05890_),
    .B(_05894_),
    .C(_05898_),
    .Y(_05899_)
  );
  NAND3X1 _13086_ (
    .A(_05889_),
    .B(_05893_),
    .C(_05897_),
    .Y(_05900_)
  );
  NAND3X1 _13087_ (
    .A(_00127_),
    .B(_05886_),
    .C(_05899_),
    .Y(_05901_)
  );
  MUX2X1 _13088_ (
    .A(_05879_),
    .B(_05878_),
    .S(_05901_),
    .Y(_05864_)
  );
  NAND2X1 _13089_ (
    .A(_00097_),
    .B(_05875_),
    .Y(_05902_)
  );
  NOR2X1 _13090_ (
    .A(_00101_),
    .B(_05902_),
    .Y(_05903_)
  );
  NAND3X1 _13091_ (
    .A(_00127_),
    .B(_05899_),
    .C(_05903_),
    .Y(_05904_)
  );
  NOR2X1 _13092_ (
    .A(_00110_),
    .B(_05904_),
    .Y(sfr_0.wdtifg_sw_clr )
  );
  NOR2X1 _13093_ (
    .A(_05878_),
    .B(_05904_),
    .Y(sfr_0.wdtifg_sw_set )
  );
  NOR2X1 _13094_ (
    .A(_00127_),
    .B(_00128_),
    .Y(_05905_)
  );
  INVX1 _13095_ (
    .A(_05905_),
    .Y(_05906_)
  );
  NAND2X1 _13096_ (
    .A(_05899_),
    .B(_05905_),
    .Y(_05907_)
  );
  AND2X1 _13097_ (
    .A(_00102_),
    .B(_05885_),
    .Y(_05908_)
  );
  NAND2X1 _13098_ (
    .A(_00102_),
    .B(_05885_),
    .Y(_05909_)
  );
  NOR3X1 _13099_ (
    .A(_05900_),
    .B(_05906_),
    .C(_05909_),
    .Y(_05910_)
  );
  NAND3X1 _13100_ (
    .A(_05899_),
    .B(_05905_),
    .C(_05908_),
    .Y(_05911_)
  );
  AND2X1 _13101_ (
    .A(1'h0),
    .B(_05910_),
    .Y(per_dout_sfr_2_)
  );
  AND2X1 _13102_ (
    .A(1'h0),
    .B(_05910_),
    .Y(per_dout_sfr_3_)
  );
  AND2X1 _13103_ (
    .A(1'h0),
    .B(_05910_),
    .Y(per_dout_sfr_4_)
  );
  AND2X1 _13104_ (
    .A(1'h0),
    .B(_05910_),
    .Y(per_dout_sfr_5_)
  );
  AND2X1 _13105_ (
    .A(1'h0),
    .B(_05910_),
    .Y(per_dout_sfr_6_)
  );
  AND2X1 _13106_ (
    .A(1'h0),
    .B(_05910_),
    .Y(per_dout_sfr_7_)
  );
  AND2X1 _13107_ (
    .A(1'h0),
    .B(_05910_),
    .Y(per_dout_sfr_9_)
  );
  AND2X1 _13108_ (
    .A(1'h0),
    .B(_05910_),
    .Y(per_dout_sfr_10_)
  );
  AND2X1 _13109_ (
    .A(1'h0),
    .B(_05910_),
    .Y(per_dout_sfr_11_)
  );
  AND2X1 _13110_ (
    .A(1'h0),
    .B(_05910_),
    .Y(per_dout_sfr_12_)
  );
  AND2X1 _13111_ (
    .A(1'h0),
    .B(_05910_),
    .Y(per_dout_sfr_13_)
  );
  NAND2X1 _13112_ (
    .A(_00101_),
    .B(_05875_),
    .Y(_05866_)
  );
  NOR2X1 _13113_ (
    .A(_00097_),
    .B(_05866_),
    .Y(_05867_)
  );
  NAND3X1 _13114_ (
    .A(_05899_),
    .B(_05905_),
    .C(_05867_),
    .Y(_05868_)
  );
  OAI21X1 _13115_ (
    .A(_05880_),
    .B(_05911_),
    .C(_05868_),
    .Y(per_dout_sfr_14_)
  );
  NOR2X1 _13116_ (
    .A(_05874_),
    .B(_05902_),
    .Y(_05869_)
  );
  NAND3X1 _13117_ (
    .A(_05899_),
    .B(_05905_),
    .C(_05869_),
    .Y(_05870_)
  );
  OAI21X1 _13118_ (
    .A(_05881_),
    .B(_05911_),
    .C(_05870_),
    .Y(per_dout_sfr_8_)
  );
  OAI21X1 _13119_ (
    .A(_05882_),
    .B(_05911_),
    .C(_05870_),
    .Y(per_dout_sfr_15_)
  );
  OAI21X1 _13120_ (
    .A(_05883_),
    .B(_05911_),
    .C(_05868_),
    .Y(per_dout_sfr_1_)
  );
  NAND2X1 _13121_ (
    .A(1'h0),
    .B(_05908_),
    .Y(_05871_)
  );
  OAI21X1 _13122_ (
    .A(_05884_),
    .B(_05902_),
    .C(_05866_),
    .Y(_05872_)
  );
  AOI21X1 _13123_ (
    .A(sfr_0.ie1_0_ ),
    .B(_05886_),
    .C(_05872_),
    .Y(_05873_)
  );
  AOI21X1 _13124_ (
    .A(_05871_),
    .B(_05873_),
    .C(_05907_),
    .Y(per_dout_sfr_0_)
  );
  DFFSR _13125_ (
    .CLK(dco_clk),
    .D(_05864_),
    .Q(sfr_0.ie1_0_ ),
    .R(_05865_),
    .S(1'h1)
  );
  INVX1 _13126_ (
    .A(_00104_),
    .Y(_05940_)
  );
  INVX1 _13127_ (
    .A(_00106_),
    .Y(_05941_)
  );
  INVX1 _13128_ (
    .A(_00108_),
    .Y(_05942_)
  );
  INVX1 _13129_ (
    .A(1'h0),
    .Y(_05943_)
  );
  INVX1 _13130_ (
    .A(_00097_),
    .Y(_05944_)
  );
  INVX1 _13131_ (
    .A(watchdog_0.wdtctl_0_ ),
    .Y(_05945_)
  );
  INVX1 _13132_ (
    .A(watchdog_0.wdtctl_1_ ),
    .Y(_05946_)
  );
  INVX1 _13133_ (
    .A(watchdog_0.wdtcnt_3_ ),
    .Y(_05947_)
  );
  INVX1 _13134_ (
    .A(watchdog_0.wdtcnt_2_ ),
    .Y(_05948_)
  );
  INVX1 _13135_ (
    .A(watchdog_0.wdtcnt_9_ ),
    .Y(_05949_)
  );
  INVX1 _13136_ (
    .A(watchdog_0.wdtcnt_10_ ),
    .Y(_05950_)
  );
  INVX1 _13137_ (
    .A(_00119_),
    .Y(_05951_)
  );
  INVX1 _13138_ (
    .A(sfr_0.wdtifg_sw_clr ),
    .Y(_05952_)
  );
  INVX1 _13139_ (
    .A(sfr_0.wdtifg_sw_set ),
    .Y(_05953_)
  );
  INVX1 _13140_ (
    .A(clock_module_0.por ),
    .Y(_05938_)
  );
  INVX1 _13141_ (
    .A(_00162_),
    .Y(_05939_)
  );
  NOR2X1 _13142_ (
    .A(_00127_),
    .B(_00128_),
    .Y(_05954_)
  );
  NOR2X1 _13143_ (
    .A(_00106_),
    .B(_00105_),
    .Y(_05955_)
  );
  NAND3X1 _13144_ (
    .A(_05942_),
    .B(_00107_),
    .C(_05955_),
    .Y(_05956_)
  );
  NOR2X1 _13145_ (
    .A(_00102_),
    .B(_00101_),
    .Y(_05957_)
  );
  NOR2X1 _13146_ (
    .A(_00103_),
    .B(_05940_),
    .Y(_05958_)
  );
  NAND2X1 _13147_ (
    .A(_05957_),
    .B(_05958_),
    .Y(_05959_)
  );
  NOR2X1 _13148_ (
    .A(_05956_),
    .B(_05959_),
    .Y(_05960_)
  );
  NAND3X1 _13149_ (
    .A(_05943_),
    .B(_00126_),
    .C(_05944_),
    .Y(_05961_)
  );
  NOR2X1 _13150_ (
    .A(_00098_),
    .B(_00109_),
    .Y(_05962_)
  );
  NOR2X1 _13151_ (
    .A(_00100_),
    .B(_00099_),
    .Y(_05963_)
  );
  NAND2X1 _13152_ (
    .A(_05962_),
    .B(_05963_),
    .Y(_05964_)
  );
  NOR2X1 _13153_ (
    .A(_05961_),
    .B(_05964_),
    .Y(_05965_)
  );
  NOR2X1 _13154_ (
    .A(_00105_),
    .B(_00108_),
    .Y(_05966_)
  );
  NOR2X1 _13155_ (
    .A(_00102_),
    .B(_05940_),
    .Y(_05967_)
  );
  OR2X1 _13156_ (
    .A(_00109_),
    .B(_00100_),
    .Y(_05968_)
  );
  NOR2X1 _13157_ (
    .A(1'h0),
    .B(_05968_),
    .Y(_05969_)
  );
  NAND3X1 _13158_ (
    .A(_05966_),
    .B(_05967_),
    .C(_05969_),
    .Y(_05970_)
  );
  NOR2X1 _13159_ (
    .A(_00101_),
    .B(_00103_),
    .Y(_05971_)
  );
  NAND3X1 _13160_ (
    .A(_05941_),
    .B(_00107_),
    .C(_05971_),
    .Y(_05972_)
  );
  NOR2X1 _13161_ (
    .A(_00098_),
    .B(_00099_),
    .Y(_05973_)
  );
  NAND3X1 _13162_ (
    .A(_00126_),
    .B(_05944_),
    .C(_05973_),
    .Y(_05974_)
  );
  OR2X1 _13163_ (
    .A(_05972_),
    .B(_05974_),
    .Y(_05975_)
  );
  NOR2X1 _13164_ (
    .A(_05970_),
    .B(_05975_),
    .Y(_05976_)
  );
  OAI21X1 _13165_ (
    .A(_00127_),
    .B(_00128_),
    .C(_05976_),
    .Y(_05977_)
  );
  MUX2X1 _13166_ (
    .A(watchdog_0.wdtctl_0_ ),
    .B(_00110_),
    .S(_05977_),
    .Y(_05978_)
  );
  INVX1 _13167_ (
    .A(_05978_),
    .Y(_05929_)
  );
  MUX2X1 _13168_ (
    .A(watchdog_0.wdtctl_1_ ),
    .B(_00117_),
    .S(_05977_),
    .Y(_05979_)
  );
  INVX1 _13169_ (
    .A(_05979_),
    .Y(_05930_)
  );
  MUX2X1 _13170_ (
    .A(watchdog_0.wdtctl_2_ ),
    .B(_00118_),
    .S(_05977_),
    .Y(_05980_)
  );
  INVX1 _13171_ (
    .A(_05980_),
    .Y(_05931_)
  );
  AND2X1 _13172_ (
    .A(watchdog_0.wdtctl_3_ ),
    .B(_05977_),
    .Y(_05932_)
  );
  MUX2X1 _13173_ (
    .A(watchdog_0.wdtctl_4_ ),
    .B(_00120_),
    .S(_05977_),
    .Y(_05981_)
  );
  INVX1 _13174_ (
    .A(_05981_),
    .Y(_05933_)
  );
  AND2X1 _13175_ (
    .A(watchdog_0.wdtctl_5_ ),
    .B(_05977_),
    .Y(_05934_)
  );
  AND2X1 _13176_ (
    .A(sfr_0.UNUSED_wdtnmies ),
    .B(_05977_),
    .Y(_05935_)
  );
  MUX2X1 _13177_ (
    .A(watchdog_0.wdtctl_7_ ),
    .B(_00123_),
    .S(_05977_),
    .Y(_05982_)
  );
  INVX1 _13178_ (
    .A(_05982_),
    .Y(_05936_)
  );
  NAND2X1 _13179_ (
    .A(watchdog_0.wdtcnt_3_ ),
    .B(watchdog_0.wdtcnt_2_ ),
    .Y(_05983_)
  );
  NAND2X1 _13180_ (
    .A(watchdog_0.wdtcnt_5_ ),
    .B(watchdog_0.wdtcnt_4_ ),
    .Y(_05984_)
  );
  NAND2X1 _13181_ (
    .A(watchdog_0.wdtcnt_0_ ),
    .B(watchdog_0.wdtcnt_1_ ),
    .Y(_05985_)
  );
  NOR3X1 _13182_ (
    .A(_05983_),
    .B(_05984_),
    .C(_05985_),
    .Y(_05986_)
  );
  AND2X1 _13183_ (
    .A(watchdog_0.wdtcnt_7_ ),
    .B(watchdog_0.wdtcnt_8_ ),
    .Y(_05987_)
  );
  NAND3X1 _13184_ (
    .A(watchdog_0.wdtcnt_6_ ),
    .B(_05986_),
    .C(_05987_),
    .Y(_05988_)
  );
  NOR2X1 _13185_ (
    .A(_05949_),
    .B(_05988_),
    .Y(_05989_)
  );
  NAND3X1 _13186_ (
    .A(watchdog_0.wdtcnt_12_ ),
    .B(watchdog_0.wdtcnt_11_ ),
    .C(watchdog_0.wdtcnt_10_ ),
    .Y(_05990_)
  );
  NOR3X1 _13187_ (
    .A(_05949_),
    .B(_05988_),
    .C(_05990_),
    .Y(_05991_)
  );
  NAND3X1 _13188_ (
    .A(watchdog_0.wdtcnt_13_ ),
    .B(watchdog_0.wdtcnt_14_ ),
    .C(_05991_),
    .Y(_05992_)
  );
  XOR2X1 _13189_ (
    .A(watchdog_0.wdtcnt_15_ ),
    .B(_05992_),
    .Y(_05993_)
  );
  XNOR2X1 _13190_ (
    .A(watchdog_0.wdtcnt_15_ ),
    .B(_05992_),
    .Y(_05994_)
  );
  NOR2X1 _13191_ (
    .A(watchdog_0.wdtctl_0_ ),
    .B(watchdog_0.wdtctl_1_ ),
    .Y(_05995_)
  );
  NAND2X1 _13192_ (
    .A(_05945_),
    .B(_05946_),
    .Y(_05996_)
  );
  XOR2X1 _13193_ (
    .A(watchdog_0.wdtcnt_13_ ),
    .B(_05991_),
    .Y(_05997_)
  );
  XNOR2X1 _13194_ (
    .A(watchdog_0.wdtcnt_13_ ),
    .B(_05991_),
    .Y(_05998_)
  );
  NAND2X1 _13195_ (
    .A(watchdog_0.wdtctl_0_ ),
    .B(watchdog_0.wdtctl_1_ ),
    .Y(_05999_)
  );
  AND2X1 _13196_ (
    .A(_05949_),
    .B(_05988_),
    .Y(_06000_)
  );
  OAI21X1 _13197_ (
    .A(_05949_),
    .B(_05988_),
    .C(watchdog_0.wdtctl_1_ ),
    .Y(_06001_)
  );
  XNOR2X1 _13198_ (
    .A(watchdog_0.wdtcnt_9_ ),
    .B(_05988_),
    .Y(_06002_)
  );
  OAI21X1 _13199_ (
    .A(watchdog_0.wdtctl_0_ ),
    .B(_06002_),
    .C(watchdog_0.wdtctl_1_ ),
    .Y(_06003_)
  );
  OAI21X1 _13200_ (
    .A(_06000_),
    .B(_06001_),
    .C(_05999_),
    .Y(_06004_)
  );
  AOI21X1 _13201_ (
    .A(watchdog_0.wdtctl_0_ ),
    .B(_05997_),
    .C(_06004_),
    .Y(_06005_)
  );
  OAI21X1 _13202_ (
    .A(_05945_),
    .B(_05998_),
    .C(_06003_),
    .Y(_06006_)
  );
  AOI21X1 _13203_ (
    .A(_05994_),
    .B(_05995_),
    .C(_06006_),
    .Y(_06007_)
  );
  OAI21X1 _13204_ (
    .A(_05993_),
    .B(_05996_),
    .C(_06005_),
    .Y(_06008_)
  );
  MUX2X1 _13205_ (
    .A(_00048_),
    .B(_00163_),
    .S(watchdog_0.wdtctl_2_ ),
    .Y(_06009_)
  );
  OR2X1 _13206_ (
    .A(watchdog_0.wdtctl_7_ ),
    .B(_00049_),
    .Y(_06010_)
  );
  NOR2X1 _13207_ (
    .A(_06009_),
    .B(_06010_),
    .Y(_06011_)
  );
  INVX1 _13208_ (
    .A(_06011_),
    .Y(_06012_)
  );
  XOR2X1 _13209_ (
    .A(watchdog_0.wdtcnt_6_ ),
    .B(_05986_),
    .Y(_06013_)
  );
  OAI21X1 _13210_ (
    .A(_05999_),
    .B(_06013_),
    .C(_06011_),
    .Y(_06014_)
  );
  INVX1 _13211_ (
    .A(_06014_),
    .Y(_06015_)
  );
  NOR2X1 _13212_ (
    .A(_00114_),
    .B(_00116_),
    .Y(_06016_)
  );
  NAND2X1 _13213_ (
    .A(_00125_),
    .B(_00112_),
    .Y(_06017_)
  );
  NOR2X1 _13214_ (
    .A(_00124_),
    .B(_00111_),
    .Y(_06018_)
  );
  NAND3X1 _13215_ (
    .A(_00113_),
    .B(_00115_),
    .C(_06018_),
    .Y(_06019_)
  );
  NOR2X1 _13216_ (
    .A(_06017_),
    .B(_06019_),
    .Y(_06020_)
  );
  AOI21X1 _13217_ (
    .A(_06016_),
    .B(_06020_),
    .C(_05977_),
    .Y(_06021_)
  );
  INVX1 _13218_ (
    .A(_06021_),
    .Y(_06022_)
  );
  AOI21X1 _13219_ (
    .A(_06008_),
    .B(_06015_),
    .C(_06021_),
    .Y(_06023_)
  );
  OAI21X1 _13220_ (
    .A(_06007_),
    .B(_06014_),
    .C(_06022_),
    .Y(_06024_)
  );
  NOR2X1 _13221_ (
    .A(_05951_),
    .B(_05977_),
    .Y(_06025_)
  );
  NAND2X1 _13222_ (
    .A(watchdog_0.wdtcnt_0_ ),
    .B(_06011_),
    .Y(_06026_)
  );
  XNOR2X1 _13223_ (
    .A(watchdog_0.wdtcnt_0_ ),
    .B(_06011_),
    .Y(_06027_)
  );
  NOR3X1 _13224_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06027_),
    .Y(_05913_)
  );
  OR2X1 _13225_ (
    .A(_05985_),
    .B(_06012_),
    .Y(_06028_)
  );
  XOR2X1 _13226_ (
    .A(watchdog_0.wdtcnt_1_ ),
    .B(_06026_),
    .Y(_06029_)
  );
  NOR3X1 _13227_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06029_),
    .Y(_05920_)
  );
  XNOR2X1 _13228_ (
    .A(_05948_),
    .B(_06028_),
    .Y(_06030_)
  );
  NOR3X1 _13229_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06030_),
    .Y(_05921_)
  );
  NOR2X1 _13230_ (
    .A(_05983_),
    .B(_06028_),
    .Y(_06031_)
  );
  OAI21X1 _13231_ (
    .A(_05948_),
    .B(_06028_),
    .C(_05947_),
    .Y(_06032_)
  );
  OAI21X1 _13232_ (
    .A(_05983_),
    .B(_06028_),
    .C(_06032_),
    .Y(_06033_)
  );
  NOR3X1 _13233_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06033_),
    .Y(_05922_)
  );
  XNOR2X1 _13234_ (
    .A(watchdog_0.wdtcnt_4_ ),
    .B(_06031_),
    .Y(_06034_)
  );
  NOR3X1 _13235_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06034_),
    .Y(_05923_)
  );
  AND2X1 _13236_ (
    .A(_05986_),
    .B(_06011_),
    .Y(_06035_)
  );
  AOI21X1 _13237_ (
    .A(watchdog_0.wdtcnt_4_ ),
    .B(_06031_),
    .C(watchdog_0.wdtcnt_5_ ),
    .Y(_06036_)
  );
  OR2X1 _13238_ (
    .A(_06035_),
    .B(_06036_),
    .Y(_06037_)
  );
  NOR3X1 _13239_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06037_),
    .Y(_05924_)
  );
  AND2X1 _13240_ (
    .A(watchdog_0.wdtcnt_6_ ),
    .B(_06035_),
    .Y(_06038_)
  );
  XNOR2X1 _13241_ (
    .A(watchdog_0.wdtcnt_6_ ),
    .B(_06035_),
    .Y(_06039_)
  );
  NOR3X1 _13242_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06039_),
    .Y(_05925_)
  );
  AND2X1 _13243_ (
    .A(watchdog_0.wdtcnt_7_ ),
    .B(_06038_),
    .Y(_06040_)
  );
  XNOR2X1 _13244_ (
    .A(watchdog_0.wdtcnt_7_ ),
    .B(_06038_),
    .Y(_06041_)
  );
  NOR3X1 _13245_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06041_),
    .Y(_05926_)
  );
  XNOR2X1 _13246_ (
    .A(watchdog_0.wdtcnt_8_ ),
    .B(_06040_),
    .Y(_06042_)
  );
  NOR3X1 _13247_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06042_),
    .Y(_05927_)
  );
  NAND2X1 _13248_ (
    .A(_05989_),
    .B(_06011_),
    .Y(_06043_)
  );
  OAI21X1 _13249_ (
    .A(_05988_),
    .B(_06012_),
    .C(_05949_),
    .Y(_06044_)
  );
  NAND2X1 _13250_ (
    .A(_06043_),
    .B(_06044_),
    .Y(_06045_)
  );
  NOR3X1 _13251_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06045_),
    .Y(_05928_)
  );
  NOR2X1 _13252_ (
    .A(_05950_),
    .B(_06043_),
    .Y(_06046_)
  );
  XNOR2X1 _13253_ (
    .A(_05950_),
    .B(_06043_),
    .Y(_06047_)
  );
  NOR3X1 _13254_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06047_),
    .Y(_05914_)
  );
  NAND2X1 _13255_ (
    .A(watchdog_0.wdtcnt_11_ ),
    .B(_06046_),
    .Y(_06048_)
  );
  XNOR2X1 _13256_ (
    .A(watchdog_0.wdtcnt_11_ ),
    .B(_06046_),
    .Y(_06049_)
  );
  NOR3X1 _13257_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06049_),
    .Y(_05915_)
  );
  XOR2X1 _13258_ (
    .A(watchdog_0.wdtcnt_12_ ),
    .B(_06048_),
    .Y(_06050_)
  );
  NOR3X1 _13259_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06050_),
    .Y(_05916_)
  );
  NAND2X1 _13260_ (
    .A(_05998_),
    .B(_06011_),
    .Y(_06051_)
  );
  OAI21X1 _13261_ (
    .A(watchdog_0.wdtcnt_13_ ),
    .B(_06011_),
    .C(_06051_),
    .Y(_06052_)
  );
  NOR3X1 _13262_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06052_),
    .Y(_05917_)
  );
  NAND3X1 _13263_ (
    .A(watchdog_0.wdtcnt_13_ ),
    .B(_05991_),
    .C(_06011_),
    .Y(_06053_)
  );
  XOR2X1 _13264_ (
    .A(watchdog_0.wdtcnt_14_ ),
    .B(_06053_),
    .Y(_06054_)
  );
  NOR3X1 _13265_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06054_),
    .Y(_05918_)
  );
  MUX2X1 _13266_ (
    .A(watchdog_0.wdtcnt_15_ ),
    .B(_05994_),
    .S(_06012_),
    .Y(_06055_)
  );
  NOR3X1 _13267_ (
    .A(_06024_),
    .B(_06025_),
    .C(_06055_),
    .Y(_05919_)
  );
  NAND2X1 _13268_ (
    .A(watchdog_0.wdtctl_4_ ),
    .B(_00084_),
    .Y(_06056_)
  );
  NAND3X1 _13269_ (
    .A(_05952_),
    .B(sfr_0.ifg1_0_ ),
    .C(_06056_),
    .Y(_06057_)
  );
  NAND3X1 _13270_ (
    .A(_05953_),
    .B(_06023_),
    .C(_06057_),
    .Y(_05937_)
  );
  NAND3X1 _13271_ (
    .A(_05954_),
    .B(_05960_),
    .C(_05965_),
    .Y(_06058_)
  );
  INVX1 _13272_ (
    .A(_06058_),
    .Y(per_dout_wdog_11_)
  );
  NAND3X1 _13273_ (
    .A(watchdog_0.wdtctl_4_ ),
    .B(sfr_0.ifg1_0_ ),
    .C(sfr_0.ie1_0_ ),
    .Y(_06059_)
  );
  INVX1 _13274_ (
    .A(_06059_),
    .Y(frontend_0.wdt_irq )
  );
  AOI22X1 _13275_ (
    .A(watchdog_0.wdtctl_4_ ),
    .B(_06022_),
    .C(_06023_),
    .D(_05953_),
    .Y(_05912_)
  );
  NOR2X1 _13276_ (
    .A(_05945_),
    .B(_06058_),
    .Y(per_dout_wdog_0_)
  );
  NOR2X1 _13277_ (
    .A(_05946_),
    .B(_06058_),
    .Y(per_dout_wdog_1_)
  );
  AND2X1 _13278_ (
    .A(watchdog_0.wdtctl_2_ ),
    .B(per_dout_wdog_11_),
    .Y(per_dout_wdog_2_)
  );
  AND2X1 _13279_ (
    .A(watchdog_0.wdtctl_3_ ),
    .B(per_dout_wdog_11_),
    .Y(per_dout_wdog_3_)
  );
  AND2X1 _13280_ (
    .A(watchdog_0.wdtctl_4_ ),
    .B(per_dout_wdog_11_),
    .Y(per_dout_wdog_4_)
  );
  AND2X1 _13281_ (
    .A(watchdog_0.wdtctl_5_ ),
    .B(per_dout_wdog_11_),
    .Y(per_dout_wdog_5_)
  );
  AND2X1 _13282_ (
    .A(sfr_0.UNUSED_wdtnmies ),
    .B(per_dout_wdog_11_),
    .Y(per_dout_wdog_6_)
  );
  AND2X1 _13283_ (
    .A(watchdog_0.wdtctl_7_ ),
    .B(per_dout_wdog_11_),
    .Y(per_dout_wdog_7_)
  );
  DFFSR _13284_ (
    .CLK(dco_clk),
    .D(_05912_),
    .Q(clock_module_0.wdt_reset ),
    .R(_05938_),
    .S(1'h1)
  );
  DFFSR _13285_ (
    .CLK(dco_clk),
    .D(_05937_),
    .Q(sfr_0.ifg1_0_ ),
    .R(_05938_),
    .S(1'h1)
  );
  DFFSR _13286_ (
    .CLK(dco_clk),
    .D(_05913_),
    .Q(watchdog_0.wdtcnt_0_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13287_ (
    .CLK(dco_clk),
    .D(_05920_),
    .Q(watchdog_0.wdtcnt_1_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13288_ (
    .CLK(dco_clk),
    .D(_05921_),
    .Q(watchdog_0.wdtcnt_2_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13289_ (
    .CLK(dco_clk),
    .D(_05922_),
    .Q(watchdog_0.wdtcnt_3_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13290_ (
    .CLK(dco_clk),
    .D(_05923_),
    .Q(watchdog_0.wdtcnt_4_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13291_ (
    .CLK(dco_clk),
    .D(_05924_),
    .Q(watchdog_0.wdtcnt_5_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13292_ (
    .CLK(dco_clk),
    .D(_05925_),
    .Q(watchdog_0.wdtcnt_6_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13293_ (
    .CLK(dco_clk),
    .D(_05926_),
    .Q(watchdog_0.wdtcnt_7_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13294_ (
    .CLK(dco_clk),
    .D(_05927_),
    .Q(watchdog_0.wdtcnt_8_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13295_ (
    .CLK(dco_clk),
    .D(_05928_),
    .Q(watchdog_0.wdtcnt_9_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13296_ (
    .CLK(dco_clk),
    .D(_05914_),
    .Q(watchdog_0.wdtcnt_10_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13297_ (
    .CLK(dco_clk),
    .D(_05915_),
    .Q(watchdog_0.wdtcnt_11_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13298_ (
    .CLK(dco_clk),
    .D(_05916_),
    .Q(watchdog_0.wdtcnt_12_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13299_ (
    .CLK(dco_clk),
    .D(_05917_),
    .Q(watchdog_0.wdtcnt_13_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13300_ (
    .CLK(dco_clk),
    .D(_05918_),
    .Q(watchdog_0.wdtcnt_14_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13301_ (
    .CLK(dco_clk),
    .D(_05919_),
    .Q(watchdog_0.wdtcnt_15_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13302_ (
    .CLK(dco_clk),
    .D(_05929_),
    .Q(watchdog_0.wdtctl_0_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13303_ (
    .CLK(dco_clk),
    .D(_05930_),
    .Q(watchdog_0.wdtctl_1_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13304_ (
    .CLK(dco_clk),
    .D(_05931_),
    .Q(watchdog_0.wdtctl_2_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13305_ (
    .CLK(dco_clk),
    .D(_05932_),
    .Q(watchdog_0.wdtctl_3_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13306_ (
    .CLK(dco_clk),
    .D(_05933_),
    .Q(watchdog_0.wdtctl_4_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13307_ (
    .CLK(dco_clk),
    .D(_05934_),
    .Q(watchdog_0.wdtctl_5_ ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13308_ (
    .CLK(dco_clk),
    .D(_05935_),
    .Q(sfr_0.UNUSED_wdtnmies ),
    .R(_05939_),
    .S(1'h1)
  );
  DFFSR _13309_ (
    .CLK(dco_clk),
    .D(_05936_),
    .Q(watchdog_0.wdtctl_7_ ),
    .R(_05939_),
    .S(1'h1)
  );
endmodule
